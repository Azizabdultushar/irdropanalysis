VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  PIN DB_Inherited_Net_Expr STRING ;
  MACRO oaTaper STRING ;
  MACRO vceLastSavedModifiedCounter INTEGER ;
END PROPERTYDEFINITIONS

MACRO ACHCONX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ACHCONX2 0 0 ;
  SIZE 7.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9746 LAYER Metal1 ;
    ANTENNADIFFAREA 5.564575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2313 LAYER Metal1 ;
      ANTENNAMAXAREACAR 17.183744 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 132.86640725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.63 0.385 6.175 0.385 6.175 0.895 6.09 0.895 6.09 1.015 6.545 1.015 6.545 1.075 6.09 1.075 6.09 1.13 5.515 1.13 5.515 1.07 6.03 1.07 6.03 0.815 6.115 0.815 6.115 0.385 5.385 0.385 5.385 0.325 6.63 0.325 ;
    END
  END CON
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0522 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.07471275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.08 0.675 0.205 1.085 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1694 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.19395 LAYER Metal1 ;
      ANTENNAMAXAREACAR 0.873421 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.81670525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.58 0.695 1.76 0.925 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0522 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.805 0.775 7.265 0.895 ;
    END
  END CI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.4 0.06 7.29 0.06 7.29 0.2 7.23 0.2 7.23 0.06 6.85 0.06 6.85 0.17 6.73 0.17 6.73 0.06 5.285 0.06 5.285 0.17 5.165 0.17 5.165 0.06 4.755 0.06 4.755 0.17 4.635 0.17 4.635 0.06 1.775 0.06 1.775 0.17 1.655 0.17 1.655 0.06 1.16 0.06 1.16 0.17 1.04 0.17 1.04 0.06 0.6 0.06 0.6 0.2 0.54 0.2 0.54 0.06 0.14 0.06 0.14 0.2 0.08 0.2 0.08 0.06 0 0.06 0 -0.06 7.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.4 1.77 0 1.77 0 1.65 0.05 1.65 0.05 1.54 0.17 1.54 0.17 1.65 0.54 1.65 0.54 1.51 0.6 1.51 0.6 1.65 1.125 1.65 1.125 1.54 1.245 1.54 1.245 1.65 1.655 1.65 1.655 1.54 1.775 1.54 1.775 1.65 4.635 1.65 4.635 1.54 4.755 1.54 4.755 1.65 5.165 1.65 5.165 1.54 5.285 1.54 5.285 1.65 6.76 1.65 6.76 1.51 6.82 1.51 6.82 1.65 7.23 1.65 7.23 1.51 7.29 1.51 7.29 1.65 7.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 7.085 0.605 6.705 0.605 6.705 1.125 7.085 1.125 7.085 1.185 6.705 1.185 6.705 1.235 6.25 1.235 6.25 1.295 6.19 1.295 6.19 1.175 6.645 1.175 6.645 0.605 6.275 0.605 6.275 0.485 6.335 0.485 6.335 0.545 7.085 0.545 ;
      POLYGON 6.015 0.71 5.93 0.71 5.93 0.89 5.7 0.89 5.7 0.97 5.415 0.97 5.415 1.13 3.27 1.13 3.27 0.97 2.65 0.97 2.65 0.91 2.73 0.91 2.73 0.49 2.67 0.49 2.67 0.43 3.54 0.43 3.54 0.49 2.79 0.49 2.79 0.91 3.33 0.91 3.33 1.07 5.355 1.07 5.355 0.91 5.64 0.91 5.64 0.83 5.87 0.83 5.87 0.59 6.015 0.59 ;
      RECT 4.9 1.23 5.84 1.29 ;
      POLYGON 5.77 0.545 5.495 0.545 5.495 0.81 5.02 0.81 5.02 0.97 4.9 0.97 4.9 0.91 4.96 0.91 4.96 0.49 4.9 0.49 4.9 0.43 5.02 0.43 5.02 0.75 5.435 0.75 5.435 0.485 5.77 0.485 ;
      POLYGON 5.335 0.65 5.12 0.65 5.12 0.33 4.8 0.33 4.8 0.49 4.21 0.49 4.21 0.91 4.27 0.91 4.27 0.97 4.15 0.97 4.15 0.43 4.74 0.43 4.74 0.27 5.18 0.27 5.18 0.59 5.335 0.59 ;
      POLYGON 4.85 0.79 4.38 0.79 4.38 0.65 4.32 0.65 4.32 0.59 4.44 0.59 4.44 0.73 4.73 0.73 4.73 0.59 4.85 0.59 ;
      POLYGON 4.535 0.33 4.05 0.33 4.05 0.97 3.79 0.97 3.79 0.91 3.99 0.91 3.99 0.33 3.155 0.33 3.155 0.27 4.535 0.27 ;
      POLYGON 4.535 1.45 1.89 1.45 1.89 1.44 0.805 1.44 0.805 0.63 0.775 0.63 0.775 0.57 0.895 0.57 0.895 0.63 0.865 0.63 0.865 1.38 1.95 1.38 1.95 1.39 4.535 1.39 ;
      POLYGON 4.145 1.29 3.11 1.29 3.11 1.13 2.21 1.13 2.21 1.095 1.97 1.095 1.97 0.695 2.14 0.695 2.14 0.43 2.26 0.43 2.26 0.49 2.2 0.49 2.2 0.755 2.03 0.755 2.03 1.035 2.27 1.035 2.27 1.07 3.17 1.07 3.17 1.23 4.145 1.23 ;
      POLYGON 3.89 0.81 3.83 0.81 3.83 0.75 3.59 0.75 3.59 0.65 3.25 0.65 3.25 0.59 3.65 0.59 3.65 0.69 3.89 0.69 ;
      POLYGON 3.55 0.91 3.43 0.91 3.43 0.81 2.95 0.81 2.95 0.65 2.89 0.65 2.89 0.59 3.01 0.59 3.01 0.75 3.49 0.75 3.49 0.85 3.55 0.85 ;
      POLYGON 3.055 0.33 1.995 0.33 1.995 0.36 1.29 0.36 1.29 1.195 2.11 1.195 2.11 1.23 3.005 1.23 3.005 1.29 2.05 1.29 2.05 1.255 1.23 1.255 1.23 0.79 0.965 0.79 0.965 0.73 1.23 0.73 1.23 0.3 1.875 0.3 1.875 0.27 3.055 0.27 ;
      POLYGON 2.55 0.935 2.13 0.935 2.13 0.855 2.47 0.855 2.47 0.56 2.55 0.56 ;
      POLYGON 2.015 0.595 1.48 0.595 1.48 1.005 1.51 1.005 1.51 1.065 1.39 1.065 1.39 1.005 1.42 1.005 1.42 0.595 1.39 0.595 1.39 0.535 2.015 0.535 ;
      POLYGON 0.705 0.79 0.365 0.79 0.365 1.285 0.305 1.285 0.305 0.595 0.275 0.595 0.275 0.535 0.395 0.535 0.395 0.595 0.365 0.595 0.365 0.73 0.705 0.73 ;
  END
END ACHCONX2

MACRO ADDFHX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFHX1 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 3.815 0.06 3.815 0.23 3.875 0.23 3.875 0.29 3.755 0.29 3.755 0.06 2.615 0.06 2.615 0.21 2.675 0.21 2.675 0.27 2.555 0.27 2.555 0.06 2.205 0.06 2.205 0.365 2.145 0.365 2.145 0.06 1.095 0.06 1.095 0.17 0.975 0.17 0.975 0.06 0.2 0.06 0.2 0.5 0.14 0.5 0.14 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.14 1.65 0.14 1.08 0.2 1.08 0.2 1.65 0.975 1.65 0.975 1.54 1.095 1.54 1.095 1.65 2.07 1.65 2.07 1.54 2.19 1.54 2.19 1.65 2.57 1.65 2.57 1.51 2.63 1.51 2.63 1.65 3.755 1.65 3.755 1.35 3.875 1.35 3.875 1.41 3.815 1.41 3.815 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.069525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.4142395 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.38 0.61 2.21 0.61 2.21 0.55 1.605 0.55 1.605 0.435 1.765 0.435 1.765 0.49 2.27 0.49 2.27 0.55 3.38 0.55 ;
    END
  END CI
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0927 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.2427185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.78 0.79 3.74 0.79 3.74 0.92 3.66 0.92 3.66 0.77 1.915 0.77 1.915 0.715 0.88 0.715 0.88 0.655 1.975 0.655 1.975 0.71 3.78 0.71 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0927 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.4142395 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.56 0.99 3.5 0.99 3.5 0.93 1.755 0.93 1.755 0.895 1.635 0.895 1.635 0.875 1.135 0.875 1.135 0.815 1.815 0.815 1.815 0.87 3.56 0.87 ;
    END
  END B
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0965 LAYER Metal1 ;
    ANTENNADIFFAREA 2.76115 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.081675 LAYER Metal1 ;
      ANTENNAMAXAREACAR 25.66880925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 189.27456375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.405 0.66 0.14 0.66 0.14 0.92 0.405 0.92 0.405 1.29 0.345 1.29 0.345 0.98 0.08 0.98 0.08 0.73 0.06 0.73 0.06 0.6 0.345 0.6 0.345 0.52 0.405 0.52 ;
    END
  END CO
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0965 LAYER Metal1 ;
    ANTENNADIFFAREA 2.76115 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.081675 LAYER Metal1 ;
      ANTENNAMAXAREACAR 25.66880925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 189.27456375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.34 0.73 4.16 0.73 4.16 1.29 4.1 1.29 4.1 0.54 4.16 0.54 4.16 0.6 4.34 0.6 ;
    END
  END S
  OBS
    LAYER Metal1 ;
      POLYGON 4 0.79 3.94 0.79 3.94 1.25 3.315 1.25 3.315 1.31 3.255 1.31 3.255 1.25 3.115 1.25 3.115 1.31 3.055 1.31 3.055 1.19 3.88 1.19 3.88 0.45 3.055 0.45 3.055 0.42 2.995 0.42 2.995 0.36 3.115 0.36 3.115 0.39 3.33 0.39 3.33 0.33 3.39 0.33 3.39 0.39 3.94 0.39 3.94 0.73 4 0.73 ;
      POLYGON 3.15 1.09 2.955 1.09 2.955 1.31 1.76 1.31 1.76 1.255 0.58 1.255 0.58 0.82 0.24 0.82 0.24 0.76 0.58 0.76 0.58 0.315 1.445 0.315 1.445 0.275 1.925 0.275 1.925 0.335 1.505 0.335 1.505 0.5 1.445 0.5 1.445 0.375 0.64 0.375 0.64 1.195 1.56 1.195 1.56 1.03 1.62 1.03 1.62 1.195 1.76 1.195 1.76 1.03 1.82 1.03 1.82 1.25 2.895 1.25 2.895 1.03 3.15 1.03 ;
      POLYGON 2.88 0.45 2.375 0.45 2.375 0.39 2.32 0.39 2.32 0.31 2.455 0.31 2.455 0.37 2.8 0.37 2.8 0.33 2.88 0.33 ;
      POLYGON 2.795 1.15 2.305 1.15 2.305 1.07 2.715 1.07 2.715 1.03 2.795 1.03 ;
      POLYGON 1.415 1.095 1.355 1.095 1.355 1.035 0.77 1.035 0.77 0.915 0.83 0.915 0.83 0.975 1.415 0.975 ;
      RECT 0.74 0.475 1.33 0.555 ;
  END
END ADDFHX1

MACRO ADDFHX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFHX2 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.29535 LAYER Metal1 ;
    ANTENNADIFFAREA 2.9812 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.140175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.3748885 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 120.8774745 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.54 0.73 4.495 0.73 4.495 1.085 4.45 1.085 4.45 1.39 4.39 1.39 4.39 1.025 4.435 1.025 4.435 0.54 4.495 0.54 4.495 0.6 4.54 0.6 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.29535 LAYER Metal1 ;
    ANTENNADIFFAREA 2.9812 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.140175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.3748885 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 120.8774745 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.34 1.29 0.28 1.29 0.28 0.73 0.26 0.73 0.26 0.6 0.28 0.6 0.28 0.54 0.34 0.54 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0927 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.44983825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.97 0.88 2.995 0.88 2.995 0.965 1.965 0.965 1.965 1.085 1.835 1.085 1.835 0.915 1.365 0.915 1.365 0.855 1.895 0.855 1.895 0.905 2.935 0.905 2.935 0.82 3.97 0.82 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0927 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.61488675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.13 0.78 4.07 0.78 4.07 0.72 2.835 0.72 2.835 0.805 2.405 0.805 2.405 0.755 1.265 0.755 1.265 0.76 1.145 0.76 1.145 0.7 1.23 0.7 1.23 0.695 2.465 0.695 2.465 0.745 2.775 0.745 2.775 0.66 3.835 0.66 3.835 0.625 3.965 0.625 3.965 0.66 4.13 0.66 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.069525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.93203875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.67 0.56 2.65 0.56 2.65 0.645 2.59 0.645 2.59 0.585 1.835 0.585 1.835 0.435 1.965 0.435 1.965 0.525 2.59 0.525 2.59 0.5 3.67 0.5 ;
    END
  END CI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.075 1.65 0.075 0.9 0.135 0.9 0.135 1.65 0.485 1.65 0.485 1.17 0.545 1.17 0.545 1.65 1.205 1.65 1.205 1.54 1.325 1.54 1.325 1.65 2.45 1.65 2.45 1.54 2.57 1.54 2.57 1.65 2.95 1.65 2.95 1.51 3.01 1.51 3.01 1.65 4.115 1.65 4.115 1.3 4.235 1.3 4.235 1.36 4.175 1.36 4.175 1.65 4.595 1.65 4.595 1 4.655 1 4.655 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 4.7 0.06 4.7 0.52 4.64 0.52 4.64 0.06 4.205 0.06 4.205 0.16 4.265 0.16 4.265 0.22 4.145 0.22 4.145 0.06 2.92 0.06 2.92 0.16 2.98 0.16 2.98 0.22 2.86 0.22 2.86 0.06 2.51 0.06 2.51 0.4 2.45 0.4 2.45 0.06 1.325 0.06 1.325 0.17 1.205 0.17 1.205 0.06 0.545 0.06 0.545 0.52 0.485 0.52 0.485 0.06 0.135 0.06 0.135 0.52 0.075 0.52 0.075 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.335 0.925 4.29 0.925 4.29 1.2 3.695 1.2 3.695 1.26 3.635 1.26 3.635 1.2 3.495 1.2 3.495 1.26 3.435 1.26 3.435 1.14 4.23 1.14 4.23 0.4 3.3 0.4 3.3 0.34 3.71 0.34 3.71 0.28 3.77 0.28 3.77 0.34 4.29 0.34 4.29 0.805 4.335 0.805 ;
      POLYGON 3.53 1.04 3.335 1.04 3.335 1.305 2.2 1.305 2.2 1.345 2.14 1.345 2.14 1.305 0.81 1.305 0.81 0.79 0.44 0.79 0.44 0.73 0.81 0.73 0.81 0.355 1.675 0.355 1.675 0.275 2.2 0.275 2.2 0.4 2.14 0.4 2.14 0.335 1.735 0.335 1.735 0.52 1.675 0.52 1.675 0.415 0.87 0.415 0.87 1.245 1.675 1.245 1.675 1.185 1.735 1.185 1.735 1.245 2.14 1.245 2.14 1.065 2.2 1.065 2.2 1.245 3.275 1.245 3.275 0.98 3.53 0.98 ;
      POLYGON 3.185 0.4 2.625 0.4 2.625 0.32 3.105 0.32 3.105 0.28 3.185 0.28 ;
      POLYGON 3.175 1.145 2.685 1.145 2.685 1.065 3.095 1.065 3.095 1.025 3.175 1.025 ;
      RECT 0.97 0.515 1.56 0.595 ;
      POLYGON 1.53 1.135 1.45 1.135 1.45 1.095 1.035 1.095 1.035 0.975 1.115 0.975 1.115 1.015 1.53 1.015 ;
  END
END ADDFHX2

MACRO ADDFHX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFHX4 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.79665 LAYER Metal1 ;
    ANTENNADIFFAREA 3.89305 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.26325 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.62355175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 79.77207975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.34 0.73 5.285 0.73 5.285 1.06 5.215 1.06 5.215 1.39 5.155 1.39 5.155 1.06 4.805 1.06 4.805 1.39 4.745 1.39 4.745 1 5.225 1 5.225 0.555 4.745 0.555 4.745 0.415 4.805 0.415 4.805 0.495 5.165 0.495 5.165 0.415 5.225 0.415 5.225 0.495 5.285 0.495 5.285 0.6 5.34 0.6 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.79665 LAYER Metal1 ;
    ANTENNADIFFAREA 3.89305 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.26325 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.62355175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 79.77207975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.82 0.66 0.34 0.66 0.34 0.92 0.82 0.92 0.82 1.295 0.76 1.295 0.76 0.98 0.4 0.98 0.4 1.295 0.34 1.295 0.34 0.98 0.28 0.98 0.28 0.73 0.26 0.73 0.26 0.6 0.34 0.6 0.34 0.52 0.4 0.52 0.4 0.6 0.76 0.6 0.76 0.52 0.82 0.52 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.102564 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.325 0.88 3.235 0.88 3.235 0.94 2.26 0.94 2.26 0.85 1.765 0.85 1.765 0.79 2.525 0.79 2.525 0.88 3.175 0.88 3.175 0.82 4.325 0.82 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.397436 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.485 0.745 4.425 0.745 4.425 0.72 3.075 0.72 3.075 0.78 2.625 0.78 2.625 0.69 1.6 0.69 1.6 0.75 1.54 0.75 1.54 0.63 2.685 0.63 2.685 0.72 3.015 0.72 3.015 0.66 4.235 0.66 4.235 0.625 4.485 0.625 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.08775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.71794875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.015 0.56 2.915 0.56 2.915 0.62 2.795 0.62 2.795 0.56 2.765 0.56 2.765 0.53 2.235 0.53 2.235 0.435 2.365 0.435 2.365 0.47 2.825 0.47 2.825 0.5 4.015 0.5 ;
    END
  END CI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 0 1.77 0 1.65 0.135 1.65 0.135 1.045 0.195 1.045 0.195 1.65 0.545 1.65 0.545 1.08 0.605 1.08 0.605 1.65 0.935 1.65 0.935 1.205 1.055 1.205 1.055 1.265 0.995 1.265 0.995 1.65 1.635 1.65 1.635 1.51 1.695 1.51 1.695 1.65 2.715 1.65 2.715 1.54 2.835 1.54 2.835 1.65 3.185 1.65 3.185 1.54 3.305 1.54 3.305 1.65 4.47 1.65 4.47 1.3 4.59 1.3 4.59 1.36 4.53 1.36 4.53 1.65 4.95 1.65 4.95 1.16 5.01 1.16 5.01 1.65 5.36 1.65 5.36 1.135 5.42 1.135 5.42 1.65 5.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5.43 0.06 5.43 0.395 5.37 0.395 5.37 0.06 5.01 0.06 5.01 0.395 4.95 0.395 4.95 0.06 4.53 0.06 4.53 0.305 4.59 0.305 4.59 0.365 4.47 0.365 4.47 0.06 3.245 0.06 3.245 0.16 3.305 0.16 3.305 0.22 3.185 0.22 3.185 0.06 2.835 0.06 2.835 0.35 2.775 0.35 2.775 0.06 1.725 0.06 1.725 0.17 1.605 0.17 1.605 0.06 1.025 0.06 1.025 0.5 0.965 0.5 0.965 0.06 0.605 0.06 0.605 0.5 0.545 0.5 0.545 0.06 0.195 0.06 0.195 0.5 0.135 0.5 0.135 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.125 0.715 4.645 0.715 4.645 1.2 4.06 1.2 4.06 1.26 4 1.26 4 1.2 3.86 1.2 3.86 1.34 3.8 1.34 3.8 1.14 4.585 1.14 4.585 0.525 4.31 0.525 4.31 0.4 3.64 0.4 3.64 0.34 4.37 0.34 4.37 0.465 4.645 0.465 4.645 0.655 5.125 0.655 ;
      POLYGON 3.865 1.04 3.7 1.04 3.7 1.28 2.465 1.28 2.465 1.34 2.405 1.34 2.405 1.28 2.135 1.28 2.135 1.32 2.075 1.32 2.075 1.23 1.21 1.23 1.21 0.82 0.44 0.82 0.44 0.76 1.21 0.76 1.21 0.29 2.075 0.29 2.075 0.25 2.525 0.25 2.525 0.37 2.465 0.37 2.465 0.31 2.135 0.31 2.135 0.45 2.075 0.45 2.075 0.35 1.27 0.35 1.27 1.17 2.075 1.17 2.075 0.95 2.135 0.95 2.135 1.22 3.64 1.22 3.64 0.98 3.865 0.98 ;
      RECT 2.95 0.32 3.54 0.4 ;
      RECT 2.95 1.04 3.54 1.12 ;
      RECT 1.37 0.45 1.96 0.53 ;
      POLYGON 1.93 1.07 1.85 1.07 1.85 1.03 1.4 1.03 1.4 0.91 1.48 0.91 1.48 0.95 1.93 0.95 ;
  END
END ADDFHX4

MACRO ADDFHXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFHXL 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.14875 LAYER Metal1 ;
    ANTENNADIFFAREA 2.6442 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.069525 LAYER Metal1 ;
      ANTENNAMAXAREACAR 30.90614875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 228.047465 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.34 0.73 4.145 0.73 4.145 1.405 4.085 1.405 4.085 0.51 4.145 0.51 4.145 0.6 4.34 0.6 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.14875 LAYER Metal1 ;
    ANTENNADIFFAREA 2.6442 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.069525 LAYER Metal1 ;
      ANTENNAMAXAREACAR 30.90614875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 228.047465 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.405 0.66 0.14 0.66 0.14 0.92 0.405 0.92 0.405 1.21 0.345 1.21 0.345 0.98 0.08 0.98 0.08 0.73 0.06 0.73 0.06 0.6 0.345 0.6 0.345 0.465 0.405 0.465 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0927 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.5598705 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.535 1.025 2.74 1.025 2.74 1.085 1.705 1.085 1.705 1.045 1.625 1.045 1.625 1.025 1.07 1.025 1.07 0.965 1.765 0.965 1.765 1.025 2.68 1.025 2.68 0.965 3.535 0.965 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0927 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.12944975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.765 0.895 3.635 0.895 3.635 0.865 2.58 0.865 2.58 0.925 1.865 0.925 1.865 0.865 0.965 0.865 0.965 0.925 0.905 0.925 0.905 0.805 1.915 0.805 1.915 0.825 1.985 0.825 1.985 0.865 2.52 0.865 2.52 0.805 3.765 0.805 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.069525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.961165 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.235 0.705 2.17 0.705 2.17 0.765 2.11 0.765 2.11 0.705 1.53 0.705 1.53 0.625 1.765 0.625 1.765 0.645 3.235 0.645 ;
    END
  END CI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.14 1.65 0.14 1.08 0.2 1.08 0.2 1.65 0.9 1.65 0.9 1.54 1.02 1.54 1.02 1.65 1.9 1.65 1.9 1.345 1.96 1.345 1.96 1.65 2.455 1.65 2.455 1.54 2.575 1.54 2.575 1.65 3.73 1.65 3.73 1.445 3.85 1.445 3.85 1.505 3.79 1.505 3.79 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 3.79 0.06 3.79 0.325 3.85 0.325 3.85 0.385 3.73 0.385 3.73 0.06 2.515 0.06 2.515 0.305 2.575 0.305 2.575 0.365 2.455 0.365 2.455 0.06 2.095 0.06 2.095 0.52 2.035 0.52 2.035 0.06 1.02 0.06 1.02 0.17 0.9 0.17 0.9 0.06 0.2 0.06 0.2 0.5 0.14 0.5 0.14 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.985 0.76 3.925 0.76 3.925 1.345 3.26 1.345 3.26 1.405 3.2 1.405 3.2 1.345 3.06 1.345 3.06 1.405 3 1.405 3 1.285 3.865 1.285 3.865 0.545 2.925 0.545 2.925 0.425 2.985 0.425 2.985 0.485 3.275 0.485 3.275 0.425 3.335 0.425 3.335 0.485 3.925 0.485 3.925 0.7 3.985 0.7 ;
      POLYGON 3.065 1.185 2.9 1.185 2.9 1.425 2.06 1.425 2.06 1.245 1.64 1.245 1.64 1.465 1.58 1.465 1.58 1.405 0.505 1.405 0.505 0.82 0.24 0.82 0.24 0.76 0.505 0.76 0.505 0.41 1.815 0.41 1.815 0.49 1.695 0.49 1.695 0.47 1.43 0.47 1.43 0.575 1.37 0.575 1.37 0.47 0.565 0.47 0.565 1.345 1.37 1.345 1.37 1.125 1.43 1.125 1.43 1.345 1.58 1.345 1.58 1.185 2.12 1.185 2.12 1.365 2.84 1.365 2.84 1.125 3.065 1.125 ;
      POLYGON 2.78 0.545 2.22 0.545 2.22 0.465 2.7 0.465 2.7 0.425 2.78 0.425 ;
      RECT 2.22 1.185 2.74 1.265 ;
      RECT 0.665 0.57 1.255 0.65 ;
      POLYGON 1.225 1.245 1.145 1.245 1.145 1.205 0.845 1.205 0.845 1.245 0.765 1.245 0.765 1.015 0.845 1.015 0.845 1.125 1.225 1.125 ;
  END
END ADDFHXL

MACRO ADDFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFX1 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.55905 LAYER Metal1 ;
    ANTENNADIFFAREA 1.826025 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0747 LAYER Metal1 ;
      ANTENNAMAXAREACAR 20.8708165 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 165.7831325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.94 1.11 2.93 1.11 2.93 1.415 2.87 1.415 2.87 1.11 2.86 1.11 2.86 0.98 2.87 0.98 2.87 0.245 2.93 0.245 2.93 0.98 2.94 0.98 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.55905 LAYER Metal1 ;
    ANTENNADIFFAREA 1.826025 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0747 LAYER Metal1 ;
      ANTENNAMAXAREACAR 20.8708165 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 165.7831325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.14 1.11 0.13 1.11 0.13 1.495 0.07 1.495 0.07 1.11 0.06 1.11 0.06 0.98 0.07 0.98 0.07 0.415 0.13 0.415 0.13 0.98 0.14 0.98 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0648 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.495 0.765 1.94 0.765 1.94 0.995 0.76 0.995 0.76 0.935 1.86 0.935 1.86 0.705 2.495 0.705 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0648 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.62037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.67 0.74 2.59 0.74 2.59 0.645 1.74 0.645 1.74 0.875 0.545 0.875 0.545 0.815 1.665 0.815 1.665 0.585 2.67 0.585 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.49382725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.41 0.525 1.57 0.525 1.57 0.755 1 0.755 1 0.695 1.435 0.695 1.435 0.6 1.46 0.6 1.46 0.465 2.41 0.465 ;
    END
  END CI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.37 0.335 1.37 0.335 1.65 0.6 1.65 0.6 1.44 0.66 1.44 0.66 1.65 1.4 1.65 1.4 1.44 1.46 1.44 1.46 1.65 1.765 1.65 1.765 1.44 1.83 1.44 1.83 1.65 2.66 1.65 2.66 1.075 2.72 1.075 2.72 1.65 3 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 0.06 2.725 0.06 2.725 0.365 2.665 0.365 2.665 0.06 1.87 0.06 1.87 0.25 1.81 0.25 1.81 0.06 1.43 0.06 1.43 0.365 1.37 0.365 1.37 0.06 0.71 0.06 0.71 0.365 0.65 0.365 0.65 0.06 0.335 0.06 0.335 0.66 0.275 0.66 0.275 0.06 0 0.06 0 -0.06 3 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.8 0.9 2.275 0.9 2.275 1.24 2.215 1.24 2.215 0.84 2.74 0.84 2.74 0.525 2.51 0.525 2.51 0.39 2.25 0.39 2.25 0.27 2.31 0.27 2.31 0.33 2.57 0.33 2.57 0.465 2.8 0.465 ;
      POLYGON 2.155 1.115 1.12 1.115 1.12 1.27 1.06 1.27 1.06 1.115 0.235 1.115 0.235 0.895 0.295 0.895 0.295 1.055 0.425 1.055 0.425 0.575 1.06 0.575 1.06 0.265 1.12 0.265 1.12 0.635 0.485 0.635 0.485 1.055 2.095 1.055 2.095 0.875 2.155 0.875 ;
      POLYGON 2.105 0.4 1.575 0.4 1.575 0.27 1.635 0.27 1.635 0.34 2.045 0.34 2.045 0.27 2.105 0.27 ;
      RECT 1.545 1.175 2.1 1.235 ;
      RECT 0.425 1.175 0.945 1.235 ;
      POLYGON 0.915 0.515 0.445 0.515 0.445 0.245 0.505 0.245 0.505 0.455 0.855 0.455 0.855 0.265 0.915 0.265 ;
  END
END ADDFX1

MACRO ADDFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFX2 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2238 LAYER Metal1 ;
    ANTENNADIFFAREA 2.658175 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1332 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.69519525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 124.27927925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.345 1.09 4.225 1.09 4.225 1.03 4.255 1.03 4.255 0.42 4.315 0.42 4.315 0.6 4.34 0.6 4.34 0.73 4.315 0.73 4.315 1.03 4.345 1.03 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2238 LAYER Metal1 ;
    ANTENNADIFFAREA 2.658175 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1332 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.69519525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 124.27927925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.335 1.31 0.275 1.31 0.275 0.85 0.14 0.85 0.14 0.92 0.06 0.92 0.06 0.79 0.275 0.79 0.275 0.54 0.335 0.54 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0648 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.17129625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.735 0.88 2.14 0.88 2.14 1.11 2.06 1.11 2.06 0.88 1.425 0.88 1.425 0.87 1.19 0.87 1.19 0.81 1.47 0.81 1.47 0.82 3.735 0.82 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0648 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 15.162037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.965 0.895 3.835 0.895 3.835 0.72 1.53 0.72 1.53 0.71 1.09 0.71 1.09 0.745 0.97 0.745 0.97 0.685 1.03 0.685 1.03 0.65 1.57 0.65 1.57 0.66 3.965 0.66 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 12.37654325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.515 0.56 1.635 0.56 1.635 0.435 1.765 0.435 1.765 0.5 3.515 0.5 ;
    END
  END CI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.02 0.13 1.02 0.13 1.65 0.45 1.65 0.45 1.22 0.57 1.22 0.57 1.28 0.51 1.28 0.51 1.65 0.92 1.65 0.92 1.51 0.98 1.51 0.98 1.65 2.12 1.65 2.12 1.51 2.18 1.51 2.18 1.65 2.575 1.65 2.575 1.54 2.695 1.54 2.695 1.65 3.88 1.65 3.88 1.3 4 1.3 4 1.36 3.94 1.36 3.94 1.65 4.46 1.65 4.46 1 4.52 1 4.52 1.65 4.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 0.06 4.52 0.06 4.52 0.4 4.46 0.4 4.46 0.06 3.97 0.06 3.97 0.4 3.91 0.4 3.91 0.06 2.78 0.06 2.78 0.16 2.84 0.16 2.84 0.22 2.72 0.22 2.72 0.06 2.205 0.06 2.205 0.31 2.265 0.31 2.265 0.37 2.145 0.37 2.145 0.06 1.195 0.06 1.195 0.17 1.075 0.17 1.075 0.06 0.54 0.06 0.54 0.52 0.48 0.52 0.48 0.06 0.13 0.06 0.13 0.52 0.07 0.52 0.07 0.06 0 0.06 0 -0.06 4.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.155 0.735 4.125 0.735 4.125 1.2 3.525 1.2 3.525 1.295 3.465 1.295 3.465 1.2 3.19 1.2 3.19 1.14 4.065 1.14 4.065 0.56 3.75 0.56 3.75 0.4 3.22 0.4 3.22 0.28 3.28 0.28 3.28 0.335 3.81 0.335 3.81 0.5 4.125 0.5 4.125 0.615 4.155 0.615 ;
      POLYGON 3.47 1.04 3.09 1.04 3.09 1.27 1.08 1.27 1.08 1.21 0.71 1.21 0.71 0.79 0.435 0.79 0.435 0.73 0.71 0.73 0.71 0.275 1.925 0.275 1.925 0.4 1.865 0.4 1.865 0.335 1.535 0.335 1.535 0.55 1.475 0.55 1.475 0.335 0.77 0.335 0.77 1.15 1.14 1.15 1.14 1.21 1.475 1.21 1.475 1.045 1.535 1.045 1.535 1.21 1.78 1.21 1.78 1.045 1.84 1.045 1.84 1.21 3.03 1.21 3.03 0.98 3.47 0.98 ;
      RECT 2.485 0.32 3.075 0.4 ;
      POLYGON 2.93 1.105 2.44 1.105 2.44 0.985 2.52 0.985 2.52 1.025 2.93 1.025 ;
      POLYGON 1.36 0.54 0.95 0.54 0.95 0.58 0.87 0.58 0.87 0.46 1.36 0.46 ;
      POLYGON 1.36 1.05 0.87 1.05 0.87 0.93 0.95 0.93 0.95 0.97 1.36 0.97 ;
  END
END ADDFX2

MACRO ADDFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFX4 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.79665 LAYER Metal1 ;
    ANTENNADIFFAREA 3.89305 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.26325 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.62355175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 79.77207975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.34 0.73 5.285 0.73 5.285 1.06 5.215 1.06 5.215 1.39 5.155 1.39 5.155 1.06 4.805 1.06 4.805 1.39 4.745 1.39 4.745 1 5.225 1 5.225 0.555 4.745 0.555 4.745 0.415 4.805 0.415 4.805 0.495 5.165 0.495 5.165 0.415 5.225 0.415 5.225 0.495 5.285 0.495 5.285 0.6 5.34 0.6 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.79665 LAYER Metal1 ;
    ANTENNADIFFAREA 3.89305 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.26325 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.62355175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 79.77207975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.82 0.66 0.34 0.66 0.34 0.92 0.82 0.92 0.82 1.295 0.76 1.295 0.76 0.98 0.4 0.98 0.4 1.295 0.34 1.295 0.34 0.98 0.28 0.98 0.28 0.73 0.26 0.73 0.26 0.6 0.34 0.6 0.34 0.52 0.4 0.52 0.4 0.6 0.76 0.6 0.76 0.52 0.82 0.52 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.102564 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.325 0.88 3.235 0.88 3.235 0.94 2.26 0.94 2.26 0.85 1.765 0.85 1.765 0.79 2.525 0.79 2.525 0.88 3.175 0.88 3.175 0.82 4.325 0.82 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.397436 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.485 0.745 4.425 0.745 4.425 0.72 3.075 0.72 3.075 0.78 2.625 0.78 2.625 0.69 1.6 0.69 1.6 0.75 1.54 0.75 1.54 0.63 2.685 0.63 2.685 0.72 3.015 0.72 3.015 0.66 4.235 0.66 4.235 0.625 4.485 0.625 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.08775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.71794875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.015 0.56 2.915 0.56 2.915 0.62 2.795 0.62 2.795 0.56 2.765 0.56 2.765 0.53 2.235 0.53 2.235 0.435 2.365 0.435 2.365 0.47 2.825 0.47 2.825 0.5 4.015 0.5 ;
    END
  END CI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 0 1.77 0 1.65 0.135 1.65 0.135 1.045 0.195 1.045 0.195 1.65 0.545 1.65 0.545 1.08 0.605 1.08 0.605 1.65 0.935 1.65 0.935 1.205 1.055 1.205 1.055 1.265 0.995 1.265 0.995 1.65 1.635 1.65 1.635 1.51 1.695 1.51 1.695 1.65 2.715 1.65 2.715 1.54 2.835 1.54 2.835 1.65 3.185 1.65 3.185 1.54 3.305 1.54 3.305 1.65 4.47 1.65 4.47 1.3 4.59 1.3 4.59 1.36 4.53 1.36 4.53 1.65 4.95 1.65 4.95 1.16 5.01 1.16 5.01 1.65 5.36 1.65 5.36 1.135 5.42 1.135 5.42 1.65 5.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5.43 0.06 5.43 0.395 5.37 0.395 5.37 0.06 5.01 0.06 5.01 0.395 4.95 0.395 4.95 0.06 4.53 0.06 4.53 0.305 4.59 0.305 4.59 0.365 4.47 0.365 4.47 0.06 3.245 0.06 3.245 0.16 3.305 0.16 3.305 0.22 3.185 0.22 3.185 0.06 2.835 0.06 2.835 0.35 2.775 0.35 2.775 0.06 1.725 0.06 1.725 0.17 1.605 0.17 1.605 0.06 1.025 0.06 1.025 0.5 0.965 0.5 0.965 0.06 0.605 0.06 0.605 0.5 0.545 0.5 0.545 0.06 0.195 0.06 0.195 0.5 0.135 0.5 0.135 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.125 0.715 4.645 0.715 4.645 1.2 4.06 1.2 4.06 1.26 4 1.26 4 1.2 3.86 1.2 3.86 1.34 3.8 1.34 3.8 1.14 4.585 1.14 4.585 0.525 4.31 0.525 4.31 0.4 3.64 0.4 3.64 0.34 4.37 0.34 4.37 0.465 4.645 0.465 4.645 0.655 5.125 0.655 ;
      POLYGON 3.865 1.04 3.7 1.04 3.7 1.28 2.465 1.28 2.465 1.34 2.405 1.34 2.405 1.28 2.135 1.28 2.135 1.32 2.075 1.32 2.075 1.23 1.21 1.23 1.21 0.82 0.44 0.82 0.44 0.76 1.21 0.76 1.21 0.29 2.075 0.29 2.075 0.25 2.525 0.25 2.525 0.37 2.465 0.37 2.465 0.31 2.135 0.31 2.135 0.45 2.075 0.45 2.075 0.35 1.27 0.35 1.27 1.17 2.075 1.17 2.075 0.95 2.135 0.95 2.135 1.22 3.64 1.22 3.64 0.98 3.865 0.98 ;
      RECT 2.95 0.32 3.54 0.4 ;
      RECT 2.95 1.04 3.54 1.12 ;
      RECT 1.37 0.45 1.96 0.53 ;
      POLYGON 1.93 1.07 1.85 1.07 1.85 1.03 1.4 1.03 1.4 0.91 1.48 0.91 1.48 0.95 1.93 0.95 ;
  END
END ADDFX4

MACRO ADDFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDFXL 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9353 LAYER Metal1 ;
    ANTENNADIFFAREA 2.131725 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXAREACAR 39.82098775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 296.54321 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.94 0.73 3.92 0.73 3.92 1.2 3.86 1.2 3.86 0.295 3.92 0.295 3.92 0.6 3.94 0.6 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9353 LAYER Metal1 ;
    ANTENNADIFFAREA 2.131725 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXAREACAR 39.82098775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 296.54321 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.375 0.54 0.14 0.54 0.14 0.86 0.375 0.86 0.375 1.045 0.315 1.045 0.315 0.92 0.06 0.92 0.06 0.79 0.08 0.79 0.08 0.48 0.315 0.48 0.315 0.285 0.375 0.285 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0648 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 12.175926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.36 0.88 2.03 0.88 2.03 0.905 1.765 0.905 1.765 1.085 1.58 1.085 1.58 0.905 1.055 0.905 1.055 0.785 1.115 0.785 1.115 0.845 1.97 0.845 1.97 0.82 3.36 0.82 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0648 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.513889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.54 1.005 3.46 1.005 3.46 0.72 1.335 0.72 1.335 0.705 1.185 0.705 1.185 0.685 0.955 0.685 0.955 0.73 0.83 0.73 0.83 0.67 0.895 0.67 0.895 0.625 1.235 0.625 1.235 0.645 1.395 0.645 1.395 0.66 3.54 0.66 ;
    END
  END A
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.98765425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.15 0.56 1.495 0.56 1.495 0.435 1.765 0.435 1.765 0.5 3.15 0.5 ;
    END
  END CI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 0 1.77 0 1.65 0.11 1.65 0.11 1.02 0.17 1.02 0.17 1.65 0.895 1.65 0.895 1.51 0.955 1.51 0.955 1.65 1.875 1.65 1.875 1.51 1.935 1.51 1.935 1.65 2.065 1.65 2.065 1.54 2.185 1.54 2.185 1.65 3.565 1.65 3.565 1.27 3.625 1.27 3.625 1.65 4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.65 0.06 3.65 0.39 3.59 0.39 3.59 0.06 2.395 0.06 2.395 0.16 2.455 0.16 2.455 0.22 2.335 0.22 2.335 0.06 1.98 0.06 1.98 0.365 1.92 0.365 1.92 0.06 1.055 0.06 1.055 0.17 0.935 0.17 0.935 0.06 0.13 0.06 0.13 0.38 0.07 0.38 0.07 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.73 1.17 2.885 1.17 2.885 1.23 2.825 1.23 2.825 1.11 3.67 1.11 3.67 0.55 3.43 0.55 3.43 0.36 2.8 0.36 2.8 0.3 3.49 0.3 3.49 0.49 3.73 0.49 ;
      POLYGON 2.725 1.38 1.535 1.38 1.535 1.245 0.54 1.245 0.54 0.7 0.3 0.7 0.3 0.76 0.24 0.76 0.24 0.64 0.54 0.64 0.54 0.275 1.625 0.275 1.625 0.335 1.395 0.335 1.395 0.545 1.335 0.545 1.335 0.335 0.6 0.335 0.6 1.185 1.335 1.185 1.335 1.05 1.395 1.05 1.395 1.185 1.595 1.185 1.595 1.32 2.665 1.32 2.665 1.04 2.555 1.04 2.555 0.98 2.725 0.98 ;
      POLYGON 2.69 0.38 2.635 0.38 2.635 0.4 2.14 0.4 2.14 0.38 2.1 0.38 2.1 0.3 2.22 0.3 2.22 0.32 2.555 0.32 2.555 0.3 2.69 0.3 ;
      POLYGON 2.565 1.22 2.05 1.22 2.05 1.045 2.13 1.045 2.13 1.14 2.565 1.14 ;
      POLYGON 1.22 0.525 0.795 0.525 0.795 0.565 0.715 0.565 0.715 0.445 1.22 0.445 ;
      RECT 0.7 1.005 1.22 1.085 ;
  END
END ADDFXL

MACRO ADDHX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHX1 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.27285 LAYER Metal1 ;
    ANTENNADIFFAREA 1.358 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0909 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.00275025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 109.6039605 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.14 0.935 2.13 0.935 2.13 1.29 2.05 1.29 2.05 0.395 2.13 0.395 2.13 0.77 2.14 0.77 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.27285 LAYER Metal1 ;
    ANTENNADIFFAREA 1.358 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0909 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.00275025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 109.6039605 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.14 1.11 0.13 1.11 0.13 1.4 0.07 1.4 0.07 1.11 0.06 1.11 0.06 0.98 0.07 0.98 0.07 0.28 0.13 0.28 0.13 0.98 0.14 0.98 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.2530865 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.645 0.885 0.565 0.885 0.565 0.92 0.435 0.92 0.435 0.765 0.645 0.765 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 17.45370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.84 1.14 0.84 1.14 0.455 0.835 0.455 0.835 0.345 0.49 0.345 0.49 0.705 0.23 0.705 0.23 0.625 0.43 0.625 0.43 0.285 0.895 0.285 0.895 0.395 1.2 0.395 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.235 1.65 0.235 1.475 0.295 1.475 0.295 1.65 0.705 1.65 0.705 1.37 0.765 1.37 0.765 1.65 1.04 1.65 1.04 1.12 1.1 1.12 1.1 1.65 1.845 1.65 1.845 1.12 1.905 1.12 1.905 1.65 2.2 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 1.905 0.06 1.905 0.64 1.845 0.64 1.845 0.06 1.05 0.06 1.05 0.285 0.99 0.285 0.99 0.06 0.365 0.06 0.365 0.535 0.245 0.535 0.245 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.99 0.79 1.595 0.79 1.595 1.24 1.535 1.24 1.535 0.535 1.595 0.535 1.595 0.73 1.99 0.73 ;
      POLYGON 1.785 0.31 1.34 0.31 1.34 1.24 1.28 1.24 1.28 0.25 1.785 0.25 ;
      POLYGON 1.69 1.44 1.16 1.44 1.16 1.03 0.895 1.03 0.895 1.195 0.835 1.195 0.835 0.535 0.895 0.535 0.895 0.97 1.22 0.97 1.22 1.38 1.415 1.38 1.415 0.845 1.4 0.845 1.4 0.725 1.475 0.725 1.475 1.38 1.69 1.38 ;
      POLYGON 0.765 1.045 0.53 1.045 0.53 1.305 0.47 1.305 0.47 1.045 0.23 1.045 0.23 0.765 0.29 0.765 0.29 0.985 0.705 0.985 0.705 0.505 0.585 0.505 0.585 0.445 0.765 0.445 ;
  END
END ADDHX1

MACRO ADDHX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHX2 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3331 LAYER Metal1 ;
    ANTENNADIFFAREA 1.951225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1494 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.9230255 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 65.993976 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.41 0.99 2.26 0.99 2.26 0.605 2.21 0.605 2.21 0.525 2.34 0.525 2.34 0.91 2.41 0.91 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3799 LAYER Metal1 ;
    ANTENNADIFFAREA 1.951225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1494 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.2362785 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 67.32931725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.115 0.865 1.115 0.865 1.035 1.06 1.035 1.06 0.635 0.77 0.635 0.77 0.555 1.14 0.555 ;
    END
  END CO
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.36 1.4 1.3 1.4 1.3 1.34 0.85 1.34 0.85 1.275 0.705 1.275 0.705 1.085 0.615 1.085 0.615 0.895 0.765 0.895 0.765 1.215 0.91 1.215 0.91 1.28 1.36 1.28 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 22.7160495 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.785 0.425 1.52 0.425 1.52 0.96 1.46 0.96 1.46 0.425 0.32 0.425 0.32 0.6 0.34 0.6 0.34 0.83 0.26 0.83 0.26 0.365 1.71 0.365 1.71 0.23 1.83 0.23 1.83 0.365 2.785 0.365 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.77 0 1.77 0 1.65 0.205 1.65 0.205 1.12 0.265 1.12 0.265 1.65 0.63 1.65 0.63 1.375 0.75 1.375 0.75 1.435 0.69 1.435 0.69 1.65 1.13 1.65 1.13 1.51 1.19 1.51 1.19 1.65 2.055 1.65 2.055 1.25 2.175 1.25 2.175 1.31 2.115 1.31 2.115 1.65 2.525 1.65 2.525 1.315 2.645 1.315 2.645 1.375 2.585 1.375 2.585 1.65 3 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 0.06 2.565 0.06 2.565 0.17 2.445 0.17 2.445 0.06 2.095 0.06 2.095 0.17 1.975 0.17 1.975 0.06 1.125 0.06 1.125 0.17 1.005 0.17 1.005 0.06 0.625 0.06 0.625 0.2 0.565 0.2 0.565 0.06 0 0.06 0 -0.06 3 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.81 0.63 2.78 0.63 2.78 1.15 2.1 1.15 2.1 0.985 1.78 0.985 1.78 0.865 1.84 0.865 1.84 0.925 2.16 0.925 2.16 1.09 2.72 1.09 2.72 0.63 2.69 0.63 2.69 0.57 2.81 0.57 ;
      POLYGON 2.16 0.825 2.1 0.825 2.1 0.765 1.68 0.765 1.68 1.145 1.62 1.145 1.62 0.545 1.755 0.545 1.755 0.605 1.68 0.605 1.68 0.705 2.16 0.705 ;
      POLYGON 1.955 1.37 1.46 1.37 1.46 1.18 1.3 1.18 1.3 0.63 1.24 0.63 1.24 0.57 1.36 0.57 1.36 1.12 1.52 1.12 1.52 1.31 1.955 1.31 ;
      POLYGON 0.925 0.855 0.865 0.855 0.865 0.795 0.5 0.795 0.5 1.15 0.38 1.15 0.38 1.09 0.44 1.09 0.44 0.99 0.1 0.99 0.1 0.54 0.16 0.54 0.16 0.93 0.44 0.93 0.44 0.735 0.925 0.735 ;
  END
END ADDHX2

MACRO ADDHX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHX4 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8982 LAYER Metal1 ;
    ANTENNADIFFAREA 3.3703 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.48957275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 47.69230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.695 1.02 3.635 1.02 3.635 0.875 3.34 0.875 3.34 0.92 3.26 0.92 3.26 0.875 3.14 0.875 3.14 1.25 3.08 1.25 3.08 0.815 3.26 0.815 3.26 0.79 3.28 0.79 3.28 0.63 3.07 0.63 3.07 0.57 3.66 0.57 3.66 0.63 3.34 0.63 3.34 0.815 3.695 0.815 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8982 LAYER Metal1 ;
    ANTENNADIFFAREA 3.3703 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.48957275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 47.69230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.5 0.64 1.34 0.64 1.34 1.07 1.5 1.07 1.5 1.13 1.28 1.13 1.28 1.01 0.91 1.01 0.91 0.95 1.26 0.95 1.26 0.64 0.8 0.64 0.8 0.52 0.86 0.52 0.86 0.58 1.44 0.58 1.44 0.51 1.5 0.51 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0747 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 22.89156625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.94 1.18 3.3 1.18 3.3 1.41 2.745 1.41 2.745 1.435 1.92 1.435 1.92 1.29 0.82 1.29 0.82 1.2 0.14 1.2 0.14 0.92 0.06 0.92 0.06 0.79 0.14 0.79 0.14 0.76 0.2 0.76 0.2 1.14 0.88 1.14 0.88 1.23 1.92 1.23 1.92 0.84 1.905 0.84 1.905 0.78 2.025 0.78 2.025 0.84 1.98 0.84 1.98 1.375 2.685 1.375 2.685 1.35 3.24 1.35 3.24 1.12 3.88 1.12 3.88 0.74 3.94 0.74 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.960396 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.855 0.68 1.6 0.68 1.6 0.41 1.34 0.41 1.34 0.42 0.7 0.42 0.7 0.66 0.54 0.66 0.54 0.8 0.46 0.8 0.46 0.6 0.64 0.6 0.64 0.36 1.28 0.36 1.28 0.35 1.66 0.35 1.66 0.62 1.855 0.62 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 1.77 0 1.77 0 1.65 0.14 1.65 0.14 1.3 0.2 1.3 0.2 1.65 0.6 1.65 0.6 1.54 0.72 1.54 0.72 1.65 1.145 1.65 1.145 1.54 1.265 1.54 1.265 1.65 1.76 1.65 1.76 1.39 1.82 1.39 1.82 1.65 2.845 1.65 2.845 1.51 2.905 1.51 2.905 1.65 3.4 1.65 3.4 1.28 3.46 1.28 3.46 1.65 3.87 1.65 3.87 1.51 3.93 1.51 3.93 1.65 4.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 0.06 3.895 0.06 3.895 0.17 3.775 0.17 3.775 0.06 3.395 0.06 3.395 0.2 3.335 0.2 3.335 0.06 2.945 0.06 2.945 0.17 2.825 0.17 2.825 0.06 1.82 0.06 1.82 0.49 1.76 0.49 1.76 0.06 1.18 0.06 1.18 0.26 1.12 0.26 1.12 0.06 0.54 0.06 0.54 0.5 0.48 0.5 0.48 0.06 0 0.06 0 -0.06 4.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.1 1.02 4.04 1.02 4.04 0.47 2.665 0.47 2.665 0.415 2.345 0.415 2.345 0.765 2.63 0.765 2.63 0.895 2.57 0.895 2.57 0.825 2.285 0.825 2.285 0.355 2.725 0.355 2.725 0.41 4.1 0.41 ;
      POLYGON 2.97 1.215 2.565 1.215 2.565 1.275 2.505 1.275 2.505 1.155 2.91 1.155 2.91 0.665 2.505 0.665 2.505 0.575 2.445 0.575 2.445 0.515 2.565 0.515 2.565 0.605 2.97 0.605 ;
      POLYGON 2.8 1.055 2.185 1.055 2.185 1.16 2.125 1.16 2.125 0.395 2.185 0.395 2.185 0.995 2.74 0.995 2.74 0.765 2.8 0.765 ;
      POLYGON 0.7 0.96 0.435 0.96 0.435 1.04 0.375 1.04 0.375 0.96 0.3 0.96 0.3 0.66 0.17 0.66 0.17 0.52 0.23 0.52 0.23 0.6 0.36 0.6 0.36 0.9 0.64 0.9 0.64 0.76 0.7 0.76 ;
  END
END ADDHX4

MACRO ADDHXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDHXL 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3132 LAYER Metal1 ;
    ANTENNADIFFAREA 1.463425 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0648 LAYER Metal1 ;
      ANTENNAMAXAREACAR 20.265432 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 156.8055555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.77 1.04 2.74 1.04 2.74 1.135 2.66 1.135 2.66 0.98 2.71 0.98 2.71 0.585 2.66 0.585 2.66 0.465 2.72 0.465 2.72 0.525 2.77 0.525 ;
    END
  END S
  PIN CO
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3613 LAYER Metal1 ;
    ANTENNADIFFAREA 1.463425 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0648 LAYER Metal1 ;
      ANTENNAMAXAREACAR 21.007716 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 160.64814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.435 0.34 1.23 ;
    END
  END CO
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.580247 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.865 0.91 0.74 0.91 0.74 1.135 0.66 1.135 0.66 0.79 0.785 0.79 0.785 0.76 0.865 0.76 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 22.22222225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.725 0.365 1.665 0.365 1.665 0.72 1.285 0.72 1.285 0.365 0.72 0.365 0.72 0.66 0.56 0.66 0.56 0.73 0.46 0.73 0.46 0.6 0.66 0.6 0.66 0.305 1.345 0.305 1.345 0.66 1.605 0.66 1.605 0.305 1.725 0.305 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 1.77 0 1.77 0 1.65 0.5 1.65 0.5 1.51 0.56 1.51 0.56 1.65 0.92 1.65 0.92 1.51 0.98 1.51 0.98 1.65 1.425 1.65 1.425 1.14 1.545 1.14 1.545 1.2 1.485 1.2 1.485 1.65 2.495 1.65 2.495 1.51 2.555 1.51 2.555 1.65 2.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 0.06 2.575 0.06 2.575 0.2 2.515 0.2 2.515 0.06 1.505 0.06 1.505 0.56 1.445 0.56 1.445 0.06 0.56 0.06 0.56 0.5 0.44 0.5 0.44 0.44 0.5 0.44 0.5 0.06 0 0.06 0 -0.06 2.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.61 0.745 2.48 0.745 2.48 1.105 2.125 1.105 2.125 1.045 2.42 1.045 2.42 0.745 2.145 0.745 2.145 0.56 2.02 0.56 2.02 0.44 2.08 0.44 2.08 0.5 2.205 0.5 2.205 0.685 2.61 0.685 ;
      POLYGON 2.415 0.34 1.92 0.34 1.92 0.525 1.825 0.525 1.825 0.82 1.865 0.82 1.865 1.135 1.805 1.135 1.805 0.88 1.765 0.88 1.765 0.465 1.86 0.465 1.86 0.28 2.415 0.28 ;
      POLYGON 2.32 0.905 2.025 0.905 2.025 1.295 1.645 1.295 1.645 1.04 1.31 1.04 1.31 1.135 1.25 1.135 1.25 0.88 1.125 0.88 1.125 0.465 1.185 0.465 1.185 0.82 1.31 0.82 1.31 0.98 1.705 0.98 1.705 1.235 1.965 1.235 1.965 0.72 1.925 0.72 1.925 0.66 2.045 0.66 2.045 0.845 2.32 0.845 ;
      POLYGON 1.025 1.295 0.44 1.295 0.44 0.95 0.5 0.95 0.5 1.235 0.965 1.235 0.965 0.525 0.82 0.525 0.82 0.465 1.025 0.465 ;
  END
END ADDHXL

MACRO AND2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X1 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3602 LAYER Metal1 ;
    ANTENNADIFFAREA 0.49995 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.31453 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 103.025641 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 0.755 0.73 0.755 0.73 1.33 0.67 1.33 0.67 0.755 0.65 0.755 0.65 0.58 0.67 0.58 0.67 0.325 0.73 0.325 0.73 0.58 0.74 0.58 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.27777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.565 1.11 0.34 1.11 0.34 0.78 0.44 0.78 0.44 0.98 0.565 0.98 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.05 0.71 0.145 0.98 ;
    END
  END B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 0.06 0.525 0.06 0.525 0.585 0.465 0.585 0.465 0.06 0 0.06 0 -0.06 0.8 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.77 0 1.77 0 1.65 0.04 1.65 0.04 1.5 0.17 1.5 0.17 1.65 0.465 1.65 0.465 1.21 0.525 1.21 0.525 1.65 0.8 1.65 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 0.59 0.855 0.53 0.855 0.53 0.715 0.27 0.715 0.27 1.21 0.315 1.21 0.315 1.33 0.255 1.33 0.255 1.27 0.21 1.27 0.21 0.605 0.12 0.605 0.12 0.465 0.18 0.465 0.18 0.545 0.27 0.545 0.27 0.645 0.59 0.645 ;
  END
END AND2X1

MACRO AND2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X2 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4539 LAYER Metal1 ;
    ANTENNADIFFAREA 0.66935 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.75897425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 64.076923 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 0.75 0.72 0.75 0.72 1.34 0.66 1.34 0.66 0.305 0.72 0.305 0.72 0.58 0.74 0.58 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.565 1.11 0.365 1.11 0.365 0.685 0.445 0.685 0.445 0.98 0.565 0.98 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.611111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.055 0.715 0.14 1.095 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.08 1.65 0.08 1.51 0.14 1.51 0.14 1.65 0.44 1.65 0.44 1.22 0.5 1.22 0.5 1.65 0.865 1.65 0.865 0.95 0.925 0.95 0.925 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.925 0.06 0.925 0.565 0.865 0.565 0.865 0.06 0.515 0.06 0.515 0.235 0.395 0.235 0.395 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.59 0.815 0.53 0.815 0.53 0.585 0.295 0.585 0.295 1.255 0.235 1.255 0.235 0.585 0.13 0.585 0.13 0.445 0.19 0.445 0.19 0.525 0.59 0.525 ;
  END
END AND2X2

MACRO AND2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X4 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.87745 LAYER Metal1 ;
    ANTENNADIFFAREA 1.11135 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.49957275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 59.897436 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.315 0.73 1.295 0.73 1.295 1.15 1.235 1.15 1.235 1.48 1.175 1.48 1.175 1.15 0.81 1.15 0.81 1.48 0.75 1.48 0.75 1.09 1.235 1.09 1.235 0.51 0.75 0.51 0.75 0.25 0.81 0.25 0.81 0.44 1.175 0.44 1.175 0.25 1.235 0.25 1.235 0.44 1.295 0.44 1.295 0.6 1.315 0.6 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.15384625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.76 0.515 1.085 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.897436 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.095 0.625 0.175 0.925 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.09 0.13 1.09 0.13 1.65 0.52 1.65 0.52 1.22 0.58 1.22 0.58 1.65 0.955 1.65 0.955 1.22 1.015 1.22 1.015 1.65 1.395 1.65 1.395 1.09 1.455 1.09 1.455 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.455 0.06 1.455 0.51 1.395 0.51 1.395 0.06 1.03 0.06 1.03 0.37 0.97 0.37 0.97 0.06 0.58 0.06 0.58 0.51 0.52 0.51 0.52 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.135 0.66 0.335 0.66 0.335 1.48 0.275 1.48 0.275 0.48 0.18 0.48 0.18 0.42 0.275 0.42 0.275 0.34 0.18 0.34 0.18 0.28 0.335 0.28 0.335 0.6 1.135 0.6 ;
  END
END AND2X4

MACRO AND2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X6 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2146 LAYER Metal1 ;
    ANTENNADIFFAREA 1.6285 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.92079775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 55.14529925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.975 1.37 1.915 1.37 1.915 0.96 1.565 0.96 1.565 1.37 1.505 1.37 1.505 0.96 1.155 0.96 1.155 1.37 1.095 1.37 1.095 0.9 1.66 0.9 1.66 0.585 1.08 0.585 1.08 0.275 1.14 0.275 1.14 0.525 1.49 0.525 1.49 0.275 1.55 0.275 1.55 0.525 1.9 0.525 1.9 0.275 1.96 0.275 1.96 0.585 1.72 0.585 1.72 0.79 1.74 0.79 1.74 0.9 1.975 0.9 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.71794875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.34 0.785 0.565 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.051282 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.82 0.755 0.76 0.755 0.76 0.685 0.185 0.685 0.185 0.78 0.125 0.78 0.125 0.705 0.06 0.705 0.06 0.625 0.82 0.625 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.98 0.13 0.98 0.13 1.65 0.48 1.65 0.48 1.13 0.54 1.13 0.54 1.65 0.89 1.65 0.89 1.13 0.95 1.13 0.95 1.65 1.3 1.65 1.3 1.06 1.36 1.06 1.36 1.65 1.71 1.65 1.71 1.06 1.77 1.06 1.77 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 1.755 0.06 1.755 0.395 1.695 0.395 1.695 0.06 1.345 0.06 1.345 0.395 1.285 0.395 1.285 0.06 0.935 0.06 0.935 0.395 0.875 0.395 0.875 0.06 0.23 0.06 0.23 0.565 0.17 0.565 0.17 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.465 0.75 0.98 0.75 0.98 1.07 0.745 1.07 0.745 1.37 0.685 1.37 0.685 1.07 0.335 1.07 0.335 1.37 0.275 1.37 0.275 1.01 0.92 1.01 0.92 0.565 0.48 0.565 0.48 0.325 0.54 0.325 0.54 0.5 0.98 0.5 0.98 0.69 1.465 0.69 ;
  END
END AND2X6

MACRO AND2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2X8 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.504775 LAYER Metal1 ;
    ANTENNADIFFAREA 1.93395 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.45549125 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 51.32561125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.42 1.425 2.36 1.425 2.36 1.045 2.01 1.045 2.01 1.425 1.95 1.425 1.95 1.045 1.6 1.045 1.6 1.425 1.54 1.425 1.54 1.045 1.19 1.045 1.19 1.425 1.13 1.425 1.13 0.98 2.06 0.98 2.06 0.66 1.075 0.66 1.075 0.275 1.135 0.275 1.135 0.595 1.485 0.595 1.485 0.275 1.545 0.275 1.545 0.595 1.895 0.595 1.895 0.275 1.955 0.275 1.955 0.595 2.305 0.595 2.305 0.275 2.365 0.275 2.365 0.66 2.14 0.66 2.14 0.845 2.12 0.845 2.12 0.98 2.42 0.98 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.17948725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.345 0.805 0.68 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 0.715 0.215 0.715 0.215 0.73 0.06 0.73 0.06 0.65 0.14 0.65 0.14 0.655 0.825 0.655 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 1.77 0 1.77 0 1.65 0.08 1.65 0.08 1.035 0.14 1.035 0.14 1.65 0.49 1.65 0.49 1.18 0.55 1.18 0.55 1.65 0.9 1.65 0.9 1.18 0.96 1.18 0.96 1.65 1.335 1.65 1.335 1.14 1.395 1.14 1.395 1.65 1.745 1.65 1.745 1.14 1.805 1.14 1.805 1.65 2.155 1.65 2.155 1.14 2.215 1.14 2.215 1.65 2.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 0.06 2.16 0.06 2.16 0.515 2.1 0.515 2.1 0.06 1.75 0.06 1.75 0.515 1.69 0.515 1.69 0.06 1.34 0.06 1.34 0.515 1.28 0.515 1.28 0.06 0.93 0.06 0.93 0.4 0.87 0.4 0.87 0.06 0.23 0.06 0.23 0.55 0.17 0.55 0.17 0.06 0 0.06 0 -0.06 2.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.92 0.83 0.945 0.83 0.945 1.12 0.755 1.12 0.755 1.425 0.695 1.425 0.695 1.12 0.345 1.12 0.345 1.425 0.285 1.425 0.285 1.06 0.885 1.06 0.885 0.565 0.49 0.565 0.49 0.31 0.55 0.31 0.55 0.5 0.945 0.5 0.945 0.77 1.92 0.77 ;
  END
END AND2X8

MACRO AND2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2XL 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3294 LAYER Metal1 ;
    ANTENNADIFFAREA 0.418125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 20.33333325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 169.72222225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.73 1.185 0.66 1.185 0.66 0.68 0.65 0.68 0.65 0.6 0.66 0.6 0.66 0.48 0.73 0.48 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.41 0.855 0.535 1.065 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.07 0.7 0.15 0.975 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.77 0 1.77 0 1.65 0.085 1.65 0.085 1.45 0.145 1.45 0.145 1.65 0.455 1.65 0.455 1.16 0.515 1.16 0.515 1.65 0.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 0.06 0.515 0.06 0.515 0.575 0.455 0.575 0.455 0.06 0 0.06 0 -0.06 0.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.58 0.765 0.31 0.765 0.31 1.185 0.25 1.185 0.25 0.6 0.14 0.6 0.14 0.48 0.2 0.48 0.2 0.54 0.31 0.54 0.31 0.705 0.58 0.705 ;
  END
END AND2XL

MACRO AND3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5341 LAYER Metal1 ;
    ANTENNADIFFAREA 0.780125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.259829 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 142.051282 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.47 1.34 1.43 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.71 0.94 1.21 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 0.98 0.52 0.98 0.52 0.87 0.34 0.87 0.34 0.92 0.26 0.92 0.26 0.79 0.6 0.79 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.16 1.17 0.06 1.17 0.06 0.98 0.08 0.98 0.08 0.69 0.16 0.69 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.435 1.65 0.435 1.51 0.495 1.51 0.495 1.65 1.04 1.65 1.04 1.31 1.1 1.31 1.1 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 1.1 0.06 1.1 0.45 1.04 0.45 1.04 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.16 0.76 1.1 0.76 1.1 0.61 0.76 0.61 0.76 1.43 0.7 1.43 0.7 1.33 0.17 1.33 0.17 1.27 0.7 1.27 0.7 0.59 0.305 0.59 0.305 0.47 0.365 0.47 0.365 0.53 0.75 0.53 0.75 0.55 1.16 0.55 ;
  END
END AND3X1

MACRO AND3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X2 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6465 LAYER Metal1 ;
    ANTENNADIFFAREA 0.8818 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.051282 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 86.5897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.73 1.32 0.73 1.32 1.42 1.26 1.42 1.26 0.66 1.145 0.66 1.145 0.48 1.205 0.48 1.205 0.6 1.34 0.6 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.965 1.085 0.915 1.085 0.915 1.455 0.835 1.455 0.835 1.005 0.965 1.005 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.575 0.735 0.495 0.735 0.495 0.64 0.34 0.64 0.34 0.73 0.26 0.73 0.26 0.56 0.575 0.56 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.16 1.04 0.06 1.04 0.06 0.79 0.08 0.79 0.08 0.56 0.16 0.56 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.44 1.65 0.44 1.3 0.5 1.3 0.5 1.65 1.015 1.65 1.015 1.3 1.075 1.3 1.075 1.65 1.465 1.65 1.465 1.03 1.525 1.03 1.525 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.41 0.06 1.41 0.46 1.35 0.46 1.35 0.06 1 0.06 1 0.46 0.94 0.46 0.94 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.045 0.73 0.735 0.73 0.735 1.325 0.675 1.325 0.675 1.2 0.325 1.2 0.325 1.295 0.205 1.295 0.205 1.235 0.265 1.235 0.265 1.14 0.675 1.14 0.675 0.46 0.28 0.46 0.28 0.34 0.34 0.34 0.34 0.4 0.735 0.4 0.735 0.67 1.045 0.67 ;
  END
END AND3X2

MACRO AND3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X4 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7914 LAYER Metal1 ;
    ANTENNADIFFAREA 1.2848 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.7641025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 56.82051275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 0.92 1.525 0.92 1.525 1.14 1.51 1.14 1.51 1.47 1.45 1.47 1.45 1.14 1.1 1.14 1.1 1.47 1.04 1.47 1.04 1.08 1.465 1.08 1.465 0.65 0.965 0.65 0.965 0.63 0.895 0.63 0.895 0.57 1.015 0.57 1.015 0.59 1.335 0.59 1.335 0.57 1.525 0.57 1.525 0.79 1.74 0.79 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 1.25 0.86 1.25 0.86 1.06 0.7 1.06 0.7 0.91 0.78 0.91 0.78 0.98 0.94 0.98 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.44 1 0.36 1 0.36 0.73 0.26 0.73 0.26 0.6 0.34 0.6 0.34 0.65 0.44 0.65 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.59 0.14 1.09 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.335 1.65 0.335 1.35 0.395 1.35 0.395 1.65 0.765 1.65 0.765 1.35 0.825 1.35 0.825 1.65 1.245 1.65 1.245 1.24 1.305 1.24 1.305 1.65 1.655 1.65 1.655 1.08 1.715 1.08 1.715 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.685 0.06 1.685 0.52 1.625 0.52 1.625 0.06 1.175 0.06 1.175 0.43 1.235 0.43 1.235 0.49 1.115 0.49 1.115 0.06 0.78 0.06 0.78 0.52 0.72 0.52 0.72 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.365 0.81 1.145 0.81 1.145 0.88 1.025 0.88 1.025 0.81 0.6 0.81 0.6 1.47 0.54 1.47 0.54 1.25 0.19 1.25 0.19 1.47 0.13 1.47 0.13 1.19 0.54 1.19 0.54 0.49 0.115 0.49 0.115 0.43 0.6 0.43 0.6 0.75 1.365 0.75 ;
  END
END AND3X4

MACRO AND3X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X6 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3559 LAYER Metal1 ;
    ANTENNADIFFAREA 1.9736 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.725926 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 60.18803425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.48 0.655 2.32 0.655 2.32 0.79 2.34 0.79 2.34 0.92 2.48 0.92 2.48 1.37 2.42 1.37 2.42 0.98 2.07 0.98 2.07 1.37 2.01 1.37 2.01 0.98 1.66 0.98 1.66 1.37 1.6 1.37 1.6 0.92 2.26 0.92 2.26 0.655 1.6 0.655 1.6 0.345 1.66 0.345 1.66 0.595 2.01 0.595 2.01 0.345 2.07 0.345 2.07 0.595 2.42 0.595 2.42 0.345 2.48 0.345 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.53 0.815 0.96 0.965 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.79487175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 0.92 1.06 0.92 1.06 0.715 0.47 0.715 0.47 0.655 1.14 0.655 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.32 0.75 1.26 0.75 1.26 0.555 0.37 0.555 0.37 0.735 0.31 0.735 0.31 0.73 0.26 0.73 0.26 0.6 0.31 0.6 0.31 0.495 1.32 0.495 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 1.77 0 1.77 0 1.65 0.165 1.65 0.165 0.98 0.225 0.98 0.225 1.65 0.575 1.65 0.575 1.25 0.635 1.25 0.635 1.65 0.985 1.65 0.985 1.25 1.045 1.25 1.045 1.65 1.395 1.65 1.395 1.25 1.455 1.25 1.455 1.65 1.805 1.65 1.805 1.08 1.865 1.08 1.865 1.65 2.215 1.65 2.215 1.08 2.275 1.08 2.275 1.65 2.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 0.06 2.275 0.06 2.275 0.465 2.215 0.465 2.215 0.06 1.865 0.06 1.865 0.465 1.805 0.465 1.805 0.06 1.455 0.06 1.455 0.17 1.335 0.17 1.335 0.06 0.265 0.06 0.265 0.335 0.325 0.335 0.325 0.395 0.205 0.395 0.205 0.06 0 0.06 0 -0.06 2.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.97 0.82 1.48 0.82 1.48 1.08 1.25 1.08 1.25 1.37 1.19 1.37 1.19 1.125 0.84 1.125 0.84 1.37 0.78 1.37 0.78 1.125 0.43 1.125 0.43 1.37 0.37 1.37 0.37 0.98 0.43 0.98 0.43 1.065 1.19 1.065 1.19 1.02 1.42 1.02 1.42 0.395 0.795 0.395 0.795 0.335 1.48 0.335 1.48 0.76 1.97 0.76 ;
  END
END AND3X6

MACRO AND3X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3X8 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.56845 LAYER Metal1 ;
    ANTENNADIFFAREA 2.241 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.72865725 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 52.35521225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.94 0.63 2.85 0.63 2.85 0.645 2.74 0.645 2.74 0.73 2.72 0.73 2.72 0.93 2.91 0.93 2.91 1.375 2.85 1.375 2.85 0.99 2.5 0.99 2.5 1.375 2.44 1.375 2.44 0.99 2.09 0.99 2.09 1.375 2.03 1.375 2.03 0.99 1.68 0.99 1.68 1.375 1.62 1.375 1.62 0.93 2.66 0.93 2.66 0.645 1.665 0.645 1.665 0.63 1.59 0.63 1.59 0.57 1.71 0.57 1.71 0.585 2 0.585 2 0.57 2.12 0.57 2.12 0.585 2.41 0.585 2.41 0.57 2.53 0.57 2.53 0.585 2.805 0.585 2.805 0.57 2.94 0.57 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.102564 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.63 0.815 0.86 0.995 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 0.92 1.06 0.92 1.06 0.715 0.58 0.715 0.58 0.655 1.14 0.655 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.76923075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.33 0.735 1.27 0.735 1.27 0.555 0.34 0.555 0.34 0.76 0.26 0.76 0.26 0.6 0.28 0.6 0.28 0.495 1.33 0.495 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.77 0 1.77 0 1.65 0.185 1.65 0.185 0.985 0.245 0.985 0.245 1.65 0.595 1.65 0.595 1.255 0.655 1.255 0.655 1.65 1.005 1.65 1.005 1.255 1.065 1.255 1.065 1.65 1.415 1.65 1.415 1.255 1.475 1.255 1.475 1.65 1.825 1.65 1.825 1.09 1.885 1.09 1.885 1.65 2.235 1.65 2.235 1.09 2.295 1.09 2.295 1.65 2.645 1.65 2.645 1.09 2.705 1.09 2.705 1.65 3 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 0.06 2.705 0.06 2.705 0.485 2.645 0.485 2.645 0.06 2.295 0.06 2.295 0.485 2.235 0.485 2.235 0.06 1.885 0.06 1.885 0.485 1.825 0.485 1.825 0.06 1.475 0.06 1.475 0.17 1.355 0.17 1.355 0.06 0.405 0.06 0.405 0.335 0.465 0.335 0.465 0.395 0.345 0.395 0.345 0.06 0 0.06 0 -0.06 3 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.39 0.805 1.49 0.805 1.49 1.08 1.27 1.08 1.27 1.375 1.21 1.375 1.21 1.155 0.86 1.155 0.86 1.375 0.8 1.375 0.8 1.155 0.45 1.155 0.45 1.375 0.39 1.375 0.39 0.985 0.45 0.985 0.45 1.095 1.21 1.095 1.21 1.02 1.43 1.02 1.43 0.395 0.815 0.395 0.815 0.335 1.49 0.335 1.49 0.745 2.39 0.745 ;
  END
END AND3X8

MACRO AND3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4911 LAYER Metal1 ;
    ANTENNADIFFAREA 0.598275 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 30.31481475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 245 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.405 1.14 1.385 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 1.12 0.86 1.12 0.86 1.06 0.72 1.06 0.72 0.76 0.8 0.76 0.8 0.98 0.94 0.98 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.46 0.91 0.34 0.91 0.34 0.98 0.26 0.98 0.26 0.79 0.38 0.79 0.38 0.6 0.46 0.6 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 1.1 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.325 1.65 0.325 1.36 0.385 1.36 0.385 1.65 0.795 1.65 0.795 1.36 0.855 1.36 0.855 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.855 0.06 0.855 0.5 0.795 0.5 0.795 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.96 0.72 0.9 0.72 0.9 0.66 0.62 0.66 0.62 1.385 0.56 1.385 0.56 1.26 0.21 1.26 0.21 1.355 0.09 1.355 0.09 1.295 0.15 1.295 0.15 1.2 0.56 1.2 0.56 0.5 0.165 0.5 0.165 0.38 0.225 0.38 0.225 0.44 0.62 0.44 0.62 0.6 0.96 0.6 ;
  END
END AND3XL

MACRO AND4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5703 LAYER Metal1 ;
    ANTENNADIFFAREA 0.793075 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.497436 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 156.6153845 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 1.345 1.155 1.345 1.155 0.27 1.215 0.27 1.215 1.17 1.34 1.17 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.68518525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.965 0.92 0.835 0.92 0.835 0.78 0.82 0.78 0.82 0.65 0.925 0.65 0.925 0.79 0.965 0.79 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.59 1.02 0.55 1.02 0.55 1.11 0.46 1.11 0.46 0.935 0.51 0.935 0.51 0.605 0.59 0.605 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.70370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.41 0.87 0.355 0.87 0.355 0.92 0.26 0.92 0.26 0.79 0.33 0.79 0.33 0.6 0.41 0.6 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.595 0.225 0.74 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.225 0.13 1.225 0.13 1.65 0.51 1.65 0.51 1.385 0.57 1.385 0.57 1.65 0.95 1.65 0.95 1.225 1.01 1.225 1.01 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 1.01 0.06 1.01 0.39 0.95 0.39 0.95 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.06 0.69 1 0.69 1 0.55 0.71 0.55 0.71 1.225 0.805 1.225 0.805 1.345 0.745 1.345 0.745 1.285 0.245 1.285 0.245 1.225 0.65 1.225 0.65 0.5 0.085 0.5 0.085 0.44 0.71 0.44 0.71 0.49 1.06 0.49 ;
  END
END AND4X1

MACRO AND4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7143 LAYER Metal1 ;
    ANTENNADIFFAREA 1.051575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.2102565 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 95.28205125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 0.73 1.46 0.73 1.46 0.875 1.365 0.875 1.365 1.335 1.305 1.335 1.305 0.815 1.4 0.815 1.4 0.415 1.305 0.415 1.305 0.295 1.365 0.295 1.365 0.355 1.46 0.355 1.46 0.6 1.54 0.6 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.115 1.06 1.115 1.06 0.92 1 0.92 1 0.675 1.08 0.675 1.08 0.775 1.14 0.775 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.6 0.74 1.1 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.5555555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.245 0.625 0.36 1.08 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.18 1.65 0.18 1.51 0.24 1.51 0.24 1.65 0.585 1.65 0.585 1.51 0.645 1.51 0.645 1.65 1.07 1.65 1.07 1.215 1.13 1.215 1.13 1.65 1.56 1.65 1.56 0.945 1.62 0.945 1.62 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.62 0.06 1.62 0.415 1.56 0.415 1.56 0.06 1.16 0.06 1.16 0.415 1.1 0.415 1.1 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.3 0.715 1.24 0.715 1.24 0.575 0.9 0.575 0.9 1.27 0.81 1.27 0.81 1.33 0.75 1.33 0.75 1.27 0.32 1.27 0.32 1.21 0.84 1.21 0.84 0.5 0.215 0.5 0.215 0.44 0.9 0.44 0.9 0.515 1.3 0.515 ;
  END
END AND4X2

MACRO AND4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X4 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9411 LAYER Metal1 ;
    ANTENNADIFFAREA 1.45555 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.04358975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 65.17948725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 0.73 1.805 0.73 1.805 1.48 1.7 1.48 1.7 1.15 1.35 1.15 1.35 1.48 1.29 1.48 1.29 1.09 1.745 1.09 1.745 0.56 1.245 0.56 1.245 0.54 1.175 0.54 1.175 0.48 1.295 0.48 1.295 0.5 1.615 0.5 1.615 0.48 1.805 0.48 1.805 0.6 1.94 0.6 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.26 1.06 1.26 1.06 1.06 1 1.06 1 0.82 1.08 0.82 1.08 0.98 1.14 0.98 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.5 0.74 1 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 1 0.48 1 0.48 0.74 0.46 0.74 0.46 0.52 0.56 0.52 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.36 0.73 0.34 0.73 0.34 0.99 0.26 0.99 0.26 0.6 0.28 0.6 0.28 0.51 0.36 0.51 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.22 1.65 0.22 1.09 0.28 1.09 0.28 1.65 0.63 1.65 0.63 1.26 0.69 1.26 0.69 1.65 1.065 1.65 1.065 1.36 1.125 1.36 1.125 1.65 1.495 1.65 1.495 1.25 1.555 1.25 1.555 1.65 1.905 1.65 1.905 1.09 1.965 1.09 1.965 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 1.965 0.06 1.965 0.43 1.905 0.43 1.905 0.06 1.455 0.06 1.455 0.34 1.515 0.34 1.515 0.4 1.395 0.4 1.395 0.06 1.06 0.06 1.06 0.43 1 0.43 1 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.645 0.72 1.425 0.72 1.425 0.88 1.305 0.88 1.305 0.72 0.9 0.72 0.9 1.48 0.84 1.48 0.84 1.16 0.485 1.16 0.485 1.48 0.425 1.48 0.425 1.1 0.84 1.1 0.84 0.4 0.235 0.4 0.235 0.34 0.9 0.34 0.9 0.66 1.645 0.66 ;
  END
END AND4X4

MACRO AND4X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X6 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5639 LAYER Metal1 ;
    ANTENNADIFFAREA 2.6403 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.911111 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 66.5128205 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.33 1.37 3.27 1.37 3.27 0.96 2.94 0.96 2.94 1.37 2.86 1.37 2.86 0.96 2.51 0.96 2.51 1.37 2.45 1.37 2.45 0.9 2.86 0.9 2.86 0.585 2.245 0.585 2.245 0.275 2.305 0.275 2.305 0.525 2.655 0.525 2.655 0.275 2.715 0.275 2.715 0.525 3.065 0.525 3.065 0.275 3.125 0.275 3.125 0.585 2.92 0.585 2.92 0.79 2.94 0.79 2.94 0.9 3.33 0.9 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.35897425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 1.11 1.92 1.11 1.92 1.185 0.395 1.185 0.395 0.82 0.455 0.82 0.455 1.125 1.86 1.125 1.86 0.82 1.94 0.82 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.76 1.025 0.66 1.025 0.66 0.895 0.555 0.895 0.555 0.835 0.66 0.835 0.66 0.79 0.74 0.79 0.74 0.965 1.7 0.965 1.7 0.845 1.76 0.845 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.051282 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.565 0.705 1.515 0.705 1.515 0.865 0.84 0.865 0.84 0.805 1.455 0.805 1.455 0.705 1.435 0.705 1.435 0.625 1.565 0.625 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.165 0.685 0.86 0.685 0.86 0.41 0.94 0.41 0.94 0.605 1.165 0.605 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 1.77 0 1.77 0 1.65 0.235 1.65 0.235 1.015 0.295 1.015 0.295 1.65 0.645 1.65 0.645 1.49 0.765 1.49 0.765 1.55 0.705 1.55 0.705 1.65 1.115 1.65 1.115 1.49 1.235 1.49 1.235 1.55 1.175 1.55 1.175 1.65 1.585 1.65 1.585 1.49 1.705 1.49 1.705 1.55 1.645 1.55 1.645 1.65 2.055 1.65 2.055 1.49 2.175 1.49 2.175 1.55 2.115 1.55 2.115 1.65 2.655 1.65 2.655 1.06 2.715 1.06 2.715 1.65 3.065 1.65 3.065 1.06 3.125 1.06 3.125 1.65 3.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 0.06 2.92 0.06 2.92 0.395 2.86 0.395 2.86 0.06 2.51 0.06 2.51 0.395 2.45 0.395 2.45 0.06 1.985 0.06 1.985 0.305 2.045 0.305 2.045 0.365 1.925 0.365 1.925 0.06 0.38 0.06 0.38 0.395 0.32 0.395 0.32 0.06 0 0.06 0 -0.06 3.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.68 0.745 2.1 0.745 2.1 1.345 1.91 1.345 1.91 1.405 1.85 1.405 1.85 1.345 1.44 1.345 1.44 1.405 1.38 1.405 1.38 1.345 0.97 1.345 0.97 1.405 0.91 1.405 0.91 1.345 0.5 1.345 0.5 1.405 0.44 1.405 0.44 1.285 2.04 1.285 2.04 0.525 1.255 0.525 1.255 0.505 1.185 0.505 1.185 0.445 1.305 0.445 1.305 0.465 2.1 0.465 2.1 0.685 2.68 0.685 ;
  END
END AND4X6

MACRO AND4X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4X8 0 0 ;
  SIZE 3.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7117 LAYER Metal1 ;
    ANTENNADIFFAREA 2.851 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.34320025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 55.66280575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.505 1.345 3.445 1.345 3.445 0.96 3.095 0.96 3.095 1.345 3.035 1.345 3.035 0.96 2.685 0.96 2.685 1.345 2.625 1.345 2.625 0.96 2.275 0.96 2.275 1.345 2.215 1.345 2.215 0.9 3.06 0.9 3.06 0.555 2.14 0.555 2.14 0.54 2.065 0.54 2.065 0.48 2.2 0.48 2.2 0.495 2.475 0.495 2.475 0.48 2.595 0.48 2.595 0.495 2.885 0.495 2.885 0.48 3.005 0.48 3.005 0.495 3.28 0.495 3.28 0.48 3.415 0.48 3.415 0.54 3.34 0.54 3.34 0.555 3.12 0.555 3.12 0.79 3.14 0.79 3.14 0.9 3.505 0.9 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.35897425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.805 1.185 0.26 1.185 0.26 0.82 0.32 0.82 0.32 1.125 1.66 1.125 1.66 0.98 1.745 0.98 1.745 0.82 1.805 0.82 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.5384615 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.645 0.88 1.56 0.88 1.56 1.025 0.46 1.025 0.46 0.895 0.42 0.895 0.42 0.835 0.46 0.835 0.46 0.79 0.54 0.79 0.54 0.965 1.5 0.965 1.5 0.76 1.645 0.76 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.30769225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.38 0.865 0.67 0.865 0.67 0.805 1.32 0.805 1.32 0.705 1.235 0.705 1.235 0.625 1.38 0.625 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.135 0.705 0.86 0.705 0.86 0.4 0.94 0.4 0.94 0.625 1.135 0.625 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 1.77 0 1.77 0 1.65 0.1 1.65 0.1 1.015 0.16 1.015 0.16 1.65 0.51 1.65 0.51 1.49 0.63 1.49 0.63 1.55 0.57 1.55 0.57 1.65 0.98 1.65 0.98 1.49 1.1 1.49 1.1 1.55 1.04 1.55 1.04 1.65 1.45 1.65 1.45 1.49 1.57 1.49 1.57 1.55 1.51 1.55 1.51 1.65 1.92 1.65 1.92 1.49 2.04 1.49 2.04 1.55 1.98 1.55 1.98 1.65 2.42 1.65 2.42 1.06 2.48 1.06 2.48 1.65 2.83 1.65 2.83 1.06 2.89 1.06 2.89 1.65 3.24 1.65 3.24 1.06 3.3 1.06 3.3 1.65 3.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 0.06 3.18 0.06 3.18 0.395 3.12 0.395 3.12 0.06 2.77 0.06 2.77 0.395 2.71 0.395 2.71 0.06 2.36 0.06 2.36 0.395 2.3 0.395 2.3 0.06 1.85 0.06 1.85 0.305 1.91 0.305 1.91 0.365 1.79 0.365 1.79 0.06 0.245 0.06 0.245 0.395 0.185 0.395 0.185 0.06 0 0.06 0 -0.06 3.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.865 0.715 1.965 0.715 1.965 1.345 1.775 1.345 1.775 1.405 1.715 1.405 1.715 1.345 1.305 1.345 1.305 1.405 1.245 1.405 1.245 1.345 0.835 1.345 0.835 1.405 0.775 1.405 0.775 1.345 0.365 1.345 0.365 1.405 0.305 1.405 0.305 1.285 1.905 1.285 1.905 0.525 1.185 0.525 1.185 0.505 1.055 0.505 1.055 0.445 1.235 0.445 1.235 0.465 1.965 0.465 1.965 0.655 2.865 0.655 ;
  END
END AND4X8

MACRO AND4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND4XL 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5472 LAYER Metal1 ;
    ANTENNADIFFAREA 0.737425 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 33.77777775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 266.4814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 1.245 1.27 1.245 1.27 0.54 1.26 0.54 1.26 0.38 1.175 0.38 1.175 0.26 1.235 0.26 1.235 0.32 1.34 0.32 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.3 1.06 1.3 1.06 1.25 1 1.25 1 0.86 1.08 0.86 1.08 1.17 1.14 1.17 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 0.92 0.72 0.92 0.72 1.12 0.64 1.12 0.64 0.64 0.74 0.64 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 0.92 0.52 0.92 0.52 1.12 0.44 1.12 0.44 0.64 0.54 0.64 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.22 0.64 0.34 1.1 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.145 1.65 0.145 1.22 0.205 1.22 0.205 1.65 0.515 1.65 0.515 1.51 0.575 1.51 0.575 1.65 1.035 1.65 1.035 1.51 1.095 1.51 1.095 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 1.03 0.06 1.03 0.38 0.97 0.38 0.97 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.16 0.6 1.1 0.6 1.1 0.54 0.9 0.54 0.9 1.28 0.81 1.28 0.81 1.34 0.75 1.34 0.75 1.28 0.32 1.28 0.32 1.22 0.84 1.22 0.84 0.54 0.275 0.54 0.275 0.375 0.215 0.375 0.215 0.315 0.335 0.315 0.335 0.48 1.16 0.48 ;
  END
END AND4XL

MACRO ANTENNA
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ANTENNA 0 0 ;
  SIZE 0.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 0.6 1.77 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 0.6 0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3439 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.39 0.34 1.27 ;
    END
  END A
END ANTENNA

MACRO AO21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6271 LAYER Metal1 ;
    ANTENNADIFFAREA 0.714625 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 21.43931625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 164.102564 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.24 1.055 1.22 1.055 1.22 1.375 1.16 1.375 1.16 0.71 1.05 0.71 1.05 0.4 1.11 0.4 1.11 0.65 1.22 0.65 1.22 0.975 1.24 0.975 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.85185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.635 0.34 0.925 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.16666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.475 0.54 0.89 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.388889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.77 0.76 1.015 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.31 1.65 0.31 1.125 0.37 1.125 0.37 1.65 0.955 1.65 0.955 1.255 1.015 1.255 1.015 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 0.905 0.06 0.905 0.52 0.845 0.52 0.845 0.06 0.245 0.06 0.245 0.52 0.185 0.52 0.185 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.965 0.82 0.9 0.82 0.9 1.155 0.815 1.155 0.815 1.215 0.755 1.215 0.755 1.095 0.84 1.095 0.84 0.68 0.64 0.68 0.64 0.425 0.7 0.425 0.7 0.62 0.9 0.62 0.9 0.7 0.965 0.7 ;
      POLYGON 0.585 1.19 0.525 1.19 0.525 1.065 0.165 1.065 0.165 1.155 0.105 1.155 0.105 1.005 0.585 1.005 ;
  END
END AO21X1

MACRO AO21X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X2 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.70675 LAYER Metal1 ;
    ANTENNADIFFAREA 0.896275 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.0811965 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 88.5641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 1.48 1.265 1.48 1.265 0.73 1.26 0.73 1.26 0.66 1.2 0.66 1.2 0.395 1.26 0.395 1.26 0.6 1.34 0.6 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.59 0.34 1.09 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.615 0.835 0.535 0.835 0.535 0.54 0.46 0.54 0.46 0.41 0.54 0.41 0.54 0.46 0.615 0.46 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.9814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 0.635 0.94 1.005 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.53 1.65 0.53 1.51 0.59 1.51 0.59 1.65 1.06 1.65 1.06 1.36 1.12 1.36 1.12 1.65 1.47 1.65 1.47 1.09 1.53 1.09 1.53 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.465 0.06 1.465 0.375 1.405 0.375 1.405 0.06 1.055 0.06 1.055 0.375 0.995 0.375 0.995 0.06 0.355 0.06 0.355 0.49 0.295 0.49 0.295 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.1 1.165 0.96 1.165 0.96 1.225 0.9 1.225 0.9 1.105 1.04 1.105 1.04 0.535 0.75 0.535 0.75 0.395 0.81 0.395 0.81 0.475 1.1 0.475 ;
      RECT 0.265 1.19 0.785 1.27 ;
  END
END AO21X2

MACRO AO21X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21X4 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.005075 LAYER Metal1 ;
    ANTENNADIFFAREA 1.309 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.5903845 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 67.4358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 0.73 1.86 0.73 1.86 0.66 1.72 0.66 1.72 1.065 1.695 1.065 1.695 1.4 1.635 1.4 1.635 1.01 1.66 1.01 1.66 0.91 1.285 0.91 1.285 1.4 1.225 1.4 1.225 0.85 1.66 0.85 1.66 0.51 1.02 0.51 1.02 0.37 1.08 0.37 1.08 0.45 1.43 0.45 1.43 0.37 1.49 0.37 1.49 0.45 1.72 0.45 1.72 0.6 1.94 0.6 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.59 0.34 1.09 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 1.09 0.46 1.09 0.46 0.79 0.48 0.79 0.48 0.61 0.56 0.61 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 1.09 0.66 1.09 0.66 0.79 0.68 0.79 0.68 0.61 0.76 0.61 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.425 1.65 0.425 1.35 0.485 1.35 0.485 1.65 1.02 1.65 1.02 1.28 1.08 1.28 1.08 1.65 1.43 1.65 1.43 1.01 1.49 1.01 1.49 1.65 1.84 1.65 1.84 1.01 1.9 1.01 1.9 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.695 0.06 1.695 0.35 1.635 0.35 1.635 0.06 1.285 0.06 1.285 0.35 1.225 0.35 1.225 0.06 0.875 0.06 0.875 0.35 0.815 0.35 0.815 0.06 0.28 0.06 0.28 0.35 0.22 0.35 0.22 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.56 0.67 0.92 0.67 0.92 1.2 0.86 1.2 0.86 0.51 0.61 0.51 0.61 0.37 0.67 0.37 0.67 0.45 0.92 0.45 0.92 0.61 1.56 0.61 ;
      POLYGON 0.69 1.47 0.63 1.47 0.63 1.25 0.28 1.25 0.28 1.47 0.22 1.47 0.22 1.19 0.69 1.19 ;
  END
END AO21X4

MACRO AO21XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO21XL 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6271 LAYER Metal1 ;
    ANTENNADIFFAREA 0.676975 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 38.7098765 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 280 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.295 0.99 1.06 0.99 1.06 0.405 1.14 0.405 1.14 0.91 1.295 0.91 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.16 1.08 0.06 1.08 0.06 0.79 0.08 0.79 0.08 0.6 0.16 0.6 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.52 0.87 0.34 0.87 0.34 0.92 0.26 0.92 0.26 0.79 0.44 0.79 0.44 0.6 0.52 0.6 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 1.19 0.66 1.19 0.66 0.81 0.62 0.81 0.62 0.73 0.74 0.73 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.32 1.65 0.32 1.36 0.38 1.36 0.38 1.65 1.04 1.65 1.04 1.285 1.1 1.285 1.1 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 0.855 0.06 0.855 0.41 0.915 0.41 0.915 0.47 0.795 0.47 0.795 0.06 0.275 0.06 0.275 0.5 0.215 0.5 0.215 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.96 0.69 0.9 0.69 0.9 1.385 0.84 1.385 0.84 0.63 0.62 0.63 0.62 0.405 0.68 0.405 0.68 0.57 0.96 0.57 ;
      POLYGON 0.615 1.37 0.48 1.37 0.48 1.26 0.205 1.26 0.205 1.355 0.085 1.355 0.085 1.275 0.125 1.275 0.125 1.18 0.56 1.18 0.56 1.29 0.615 1.29 ;
  END
END AO21XL

MACRO AO22X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X1 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7252 LAYER Metal1 ;
    ANTENNADIFFAREA 0.85985 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 24.7931625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 189.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 1.3 1.345 1.3 1.345 1.44 1.285 1.44 1.285 1.3 1.235 1.3 1.235 1.17 1.285 1.17 1.285 0.275 1.345 0.275 1.345 1.17 1.365 1.17 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.9814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.41 0.945 0.81 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 12.12962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.205 0.72 0.14 0.72 0.14 1.11 0.06 1.11 0.06 0.6 0.205 0.6 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.4074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.605 0.855 0.525 0.855 0.525 0.745 0.46 0.745 0.46 0.6 0.605 0.6 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.388889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.41 0.985 0.33 0.985 0.33 0.92 0.26 0.92 0.26 0.79 0.41 0.79 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.305 1.65 0.305 1.51 0.365 1.51 0.365 1.65 1.08 1.65 1.08 1.05 1.14 1.05 1.14 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.14 0.06 1.14 0.535 1.08 0.535 1.08 0.06 0.22 0.06 0.22 0.51 0.16 0.51 0.16 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.225 0.95 0.765 0.95 0.765 1.235 0.645 1.235 0.645 1.175 0.705 1.175 0.705 0.505 0.44 0.505 0.44 0.445 0.765 0.445 0.765 0.89 1.225 0.89 ;
      POLYGON 0.94 1.395 0.47 1.395 0.47 1.28 0.04 1.28 0.04 1.22 0.53 1.22 0.53 1.335 0.88 1.335 0.88 1.22 0.94 1.22 ;
  END
END AO22X1

MACRO AO22X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7356 LAYER Metal1 ;
    ANTENNADIFFAREA 1.0615 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.574359 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 98.3846155 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 1.48 1.465 1.48 1.465 1.11 1.46 1.11 1.46 0.415 1.52 0.415 1.52 0.98 1.54 0.98 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.12 1.025 1.12 1.025 0.655 1.105 0.655 1.105 0.955 1.14 0.955 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.16 1.11 0.06 1.11 0.06 0.955 0.08 0.955 0.08 0.63 0.16 0.63 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.765 1.055 0.685 1.055 0.685 0.705 0.635 0.705 0.635 0.605 0.765 0.605 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.535 1.07 0.455 1.07 0.455 0.895 0.34 0.895 0.34 0.92 0.26 0.92 0.26 0.79 0.34 0.79 0.34 0.815 0.535 0.815 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.305 1.65 0.305 1.51 0.365 1.51 0.365 1.65 1.23 1.65 1.23 1.39 1.35 1.39 1.35 1.45 1.29 1.45 1.29 1.65 1.67 1.65 1.67 1.09 1.73 1.09 1.73 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.725 0.06 1.725 0.395 1.665 0.395 1.665 0.06 1.315 0.06 1.315 0.395 1.255 0.395 1.255 0.06 0.29 0.06 0.29 0.51 0.23 0.51 0.23 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.36 0.695 1.3 0.695 1.3 0.555 0.925 0.555 0.925 1.215 0.8 1.215 0.8 1.155 0.865 1.155 0.865 0.505 0.6 0.505 0.6 0.445 0.925 0.445 0.925 0.495 1.36 0.495 ;
      POLYGON 1.095 1.375 0.54 1.375 0.54 1.28 0.04 1.28 0.04 1.22 0.6 1.22 0.6 1.315 1.035 1.315 1.035 1.22 1.095 1.22 ;
  END
END AO22X2

MACRO AO22X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22X4 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0641 LAYER Metal1 ;
    ANTENNADIFFAREA 1.5177 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.09487175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 70.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 0.73 1.92 0.73 1.92 1.305 1.86 1.305 1.86 0.975 1.51 0.975 1.51 1.305 1.45 1.305 1.45 0.915 1.86 0.915 1.86 0.55 1.315 0.55 1.315 0.53 1.245 0.53 1.245 0.47 1.365 0.47 1.365 0.49 1.685 0.49 1.685 0.47 1.805 0.47 1.805 0.49 1.92 0.49 1.92 0.6 1.94 0.6 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.31 1.085 1.035 1.085 1.035 0.895 1 0.895 1 0.815 1.12 0.815 1.12 1.005 1.31 1.005 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.52 0.34 1.02 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.52 0.74 1.02 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 1 0.46 1 0.46 0.79 0.48 0.79 0.48 0.52 0.56 0.52 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.425 1.65 0.425 1.28 0.485 1.28 0.485 1.65 1.215 1.65 1.215 1.51 1.275 1.51 1.275 1.65 1.655 1.65 1.655 1.075 1.715 1.075 1.715 1.65 2.065 1.65 2.065 0.915 2.125 0.915 2.125 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 1.965 0.06 1.965 0.33 2.025 0.33 2.025 0.39 1.905 0.39 1.905 0.06 1.525 0.06 1.525 0.33 1.585 0.33 1.585 0.39 1.465 0.39 1.465 0.06 1.105 0.06 1.105 0.42 1.045 0.42 1.045 0.06 0.28 0.06 0.28 0.42 0.22 0.42 0.22 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.74 0.715 0.9 0.715 0.9 1.24 0.84 1.24 0.84 0.42 0.6 0.42 0.6 0.36 0.9 0.36 0.9 0.655 1.74 0.655 ;
      POLYGON 1.105 1.4 0.63 1.4 0.63 1.18 0.28 1.18 0.28 1.4 0.22 1.4 0.22 1.12 0.69 1.12 0.69 1.34 1.045 1.34 1.045 1.28 1.105 1.28 ;
  END
END AO22X4

MACRO AO22XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AO22XL 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6486 LAYER Metal1 ;
    ANTENNADIFFAREA 0.76475 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 40.037037 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 310.83333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.51 0.99 1.26 0.99 1.26 0.68 1.25 0.68 1.25 0.405 1.33 0.405 1.33 0.6 1.34 0.6 1.34 0.91 1.51 0.91 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.23 1.06 1.23 1.06 0.87 1 0.87 1 0.79 1.14 0.79 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 1.1 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.595 0.74 1.095 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.23 0.54 0.73 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.41 1.65 0.41 1.36 0.47 1.36 0.47 1.65 1.255 1.65 1.255 1.33 1.315 1.33 1.315 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.075 0.06 1.075 0.41 1.135 0.41 1.135 0.47 1.015 0.47 1.015 0.06 0.265 0.06 0.265 0.5 0.205 0.5 0.205 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.145 0.69 0.9 0.69 0.9 1.385 0.84 1.385 0.84 0.495 0.64 0.495 0.64 0.435 0.9 0.435 0.9 0.63 1.085 0.63 1.085 0.57 1.145 0.57 ;
      POLYGON 1.135 1.45 1.06 1.45 1.06 1.545 0.615 1.545 0.615 1.26 0.295 1.26 0.295 1.355 0.175 1.355 0.175 1.295 0.235 1.295 0.235 1.2 0.675 1.2 0.675 1.485 1 1.485 1 1.39 1.135 1.39 ;
  END
END AO22XL

MACRO AOI211X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5721 LAYER Metal1 ;
    ANTENNADIFFAREA 0.817 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.3 1.18 1.095 1.18 1.095 1.48 1.035 1.48 1.035 1.12 1.24 1.12 1.24 0.54 0.63 0.54 0.63 0.5 0.58 0.5 0.58 0.44 0.7 0.44 0.7 0.48 1.06 0.48 1.06 0.41 1.14 0.41 1.14 0.48 1.3 0.48 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 1.1 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.6 0.54 1.1 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.84 0.72 0.74 0.72 0.74 1.04 0.66 1.04 0.66 0.64 0.84 0.64 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.02 1.06 1.02 1.06 0.87 0.94 0.87 0.94 0.64 1.02 0.64 1.02 0.79 1.14 0.79 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.45 1.65 0.45 1.36 0.51 1.36 0.51 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 0.86 0.06 0.86 0.32 0.92 0.32 0.92 0.38 0.8 0.38 0.8 0.06 0.305 0.06 0.305 0.41 0.245 0.41 0.245 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.715 1.48 0.655 1.48 0.655 1.26 0.305 1.26 0.305 1.48 0.245 1.48 0.245 1.2 0.715 1.2 ;
  END
END AOI211X1

MACRO AOI211X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9703 LAYER Metal1 ;
    ANTENNADIFFAREA 1.43645 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.755 0.505 1.685 0.505 1.685 0.525 1.14 0.525 1.14 0.945 1.725 0.945 1.725 1.225 1.665 1.225 1.665 1.005 1.08 1.005 1.08 0.73 1.06 0.73 1.06 0.525 0.62 0.525 0.62 0.505 0.55 0.505 0.55 0.445 0.67 0.445 0.67 0.465 1.195 0.465 1.195 0.445 1.315 0.445 1.315 0.465 1.635 0.465 1.635 0.445 1.755 0.445 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.4615385 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.525 0.805 0.895 0.915 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.84615375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.625 0.905 0.705 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.845 1.435 0.845 1.435 0.705 1.24 0.705 1.24 0.625 1.6 0.625 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.7 0.625 1.965 0.795 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.995 0.13 0.995 0.13 1.65 0.48 1.65 0.48 1.265 0.54 1.265 0.54 1.65 0.92 1.65 0.92 1.51 0.98 1.51 0.98 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.93 0.06 1.93 0.395 1.87 0.395 1.87 0.06 1.475 0.06 1.475 0.305 1.535 0.305 1.535 0.365 1.415 0.365 1.415 0.06 0.92 0.06 0.92 0.305 0.98 0.305 0.98 0.365 0.86 0.365 0.86 0.06 0.32 0.06 0.32 0.395 0.26 0.395 0.26 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.93 1.385 1.095 1.385 1.095 1.325 1.02 1.325 1.02 1.265 1.155 1.265 1.155 1.325 1.46 1.325 1.46 1.235 1.52 1.235 1.52 1.325 1.87 1.325 1.87 0.965 1.93 0.965 ;
      POLYGON 1.315 1.225 1.255 1.225 1.255 1.165 0.745 1.165 0.745 1.385 0.685 1.385 0.685 1.165 0.335 1.165 0.335 1.385 0.275 1.385 0.275 1.105 1.315 1.105 ;
  END
END AOI211X2

MACRO AOI211X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211X4 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8385 LAYER Metal1 ;
    ANTENNADIFFAREA 2.64575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.455 1.275 3.395 1.275 3.395 1.105 3.045 1.105 3.045 1.275 2.985 1.275 2.985 1.055 1.905 1.055 1.905 0.705 1.835 0.705 1.835 0.625 1.905 0.625 1.905 0.525 0.83 0.525 0.83 0.505 0.76 0.505 0.76 0.445 0.88 0.445 0.88 0.465 1.38 0.465 1.38 0.445 1.5 0.445 1.5 0.465 1.935 0.465 1.935 0.445 2.055 0.445 2.055 0.465 2.415 0.465 2.415 0.445 2.535 0.445 2.535 0.465 2.855 0.465 2.855 0.445 2.975 0.445 2.975 0.465 3.295 0.465 3.295 0.445 3.415 0.445 3.415 0.505 3.345 0.505 3.345 0.525 1.965 0.525 1.965 0.995 3.045 0.995 3.045 1.045 3.455 1.045 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.102564 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 0.815 1.425 0.895 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.065 0.815 2.565 0.895 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.365 0.825 3.285 0.825 3.285 0.705 2.985 0.705 2.985 0.625 3.365 0.625 ;
    END
  END C0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.0641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.735 0.705 0.23 0.705 0.23 0.645 0.235 0.645 0.235 0.625 0.365 0.625 0.365 0.645 1.735 0.645 ;
    END
  END A0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 1.77 0 1.77 0 1.65 0.13 1.65 0.13 1.045 0.19 1.045 0.19 1.65 0.54 1.65 0.54 1.315 0.6 1.315 0.6 1.65 0.95 1.65 0.95 1.315 1.01 1.315 1.01 1.65 1.36 1.65 1.36 1.315 1.42 1.315 1.42 1.65 1.8 1.65 1.8 1.51 1.86 1.51 1.86 1.65 3.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 0.06 3.59 0.06 3.59 0.395 3.53 0.395 3.53 0.06 3.135 0.06 3.135 0.305 3.195 0.305 3.195 0.365 3.075 0.365 3.075 0.06 2.695 0.06 2.695 0.305 2.755 0.305 2.755 0.365 2.635 0.365 2.635 0.06 2.215 0.06 2.215 0.305 2.275 0.305 2.275 0.365 2.155 0.365 2.155 0.06 1.75 0.06 1.75 0.305 1.81 0.305 1.81 0.365 1.69 0.365 1.69 0.06 1.13 0.06 1.13 0.305 1.19 0.305 1.19 0.365 1.07 0.365 1.07 0.06 0.54 0.06 0.54 0.395 0.48 0.395 0.48 0.06 0 0.06 0 -0.06 3.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.66 1.435 2.005 1.435 2.005 1.4 1.93 1.4 1.93 1.34 2.065 1.34 2.065 1.375 2.37 1.375 2.37 1.315 2.43 1.315 2.43 1.375 2.78 1.375 2.78 1.155 2.84 1.155 2.84 1.375 3.19 1.375 3.19 1.205 3.25 1.205 3.25 1.375 3.6 1.375 3.6 1.045 3.66 1.045 ;
      POLYGON 2.635 1.275 2.575 1.275 2.575 1.215 2.225 1.215 2.225 1.275 2.165 1.275 2.165 1.215 1.625 1.215 1.625 1.435 1.565 1.435 1.565 1.215 1.215 1.215 1.215 1.435 1.155 1.435 1.155 1.215 0.805 1.215 0.805 1.435 0.745 1.435 0.745 1.215 0.395 1.215 0.395 1.435 0.335 1.435 0.335 1.155 2.635 1.155 ;
  END
END AOI211X4

MACRO AOI211XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.528875 LAYER Metal1 ;
    ANTENNADIFFAREA 0.589525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.295 1.06 1.295 1.06 0.98 1.08 0.98 1.08 0.51 0.595 0.51 0.595 0.285 0.655 0.285 0.655 0.45 1.005 0.45 1.005 0.285 1.14 0.285 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.16 0.99 0.08 0.99 0.08 0.73 0.06 0.73 0.06 0.51 0.16 0.51 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.46 0.705 0.34 0.705 0.34 0.99 0.26 0.99 0.26 0.61 0.46 0.61 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 0.69 0.74 0.69 0.74 0.99 0.66 0.99 0.66 0.69 0.56 0.69 0.56 0.61 0.76 0.61 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.61 0.94 1.11 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.305 1.65 0.305 1.27 0.365 1.27 0.365 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.83 0.06 0.83 0.29 0.89 0.29 0.89 0.35 0.77 0.35 0.77 0.06 0.26 0.06 0.26 0.38 0.2 0.38 0.2 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.6 1.29 0.465 1.29 0.465 1.17 0.19 1.17 0.19 1.265 0.07 1.265 0.07 1.185 0.11 1.185 0.11 1.09 0.545 1.09 0.545 1.21 0.6 1.21 ;
  END
END AOI211XL

MACRO AOI21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X1 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4656 LAYER Metal1 ;
    ANTENNADIFFAREA 0.63925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.78 1.11 0.76 1.11 0.76 1.44 0.7 1.44 0.7 1.11 0.66 1.11 0.66 0.98 0.7 0.98 0.7 0.48 0.38 0.48 0.38 0.23 0.44 0.23 0.44 0.42 0.76 0.42 0.76 0.98 0.78 0.98 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.69230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.44 0.18 0.68 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.897436 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.58 0.38 0.84 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.076923 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 0.66 0.54 0.66 0.54 0.935 0.46 0.935 0.46 0.58 0.6 0.58 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.2 0.335 1.2 0.335 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.645 0.06 0.645 0.35 0.585 0.35 0.585 0.06 0.13 0.06 0.13 0.35 0.07 0.35 0.07 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.54 1.44 0.48 1.44 0.48 1.14 0.13 1.14 0.13 1.44 0.07 1.44 0.07 1.08 0.54 1.08 ;
  END
END AOI21X1

MACRO AOI21X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X2 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.345 0.06 1.345 0.36 1.285 0.36 1.285 0.06 0.9 0.06 0.9 0.27 0.96 0.27 0.96 0.33 0.84 0.33 0.84 0.06 0.285 0.06 0.285 0.36 0.225 0.36 0.225 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.33 1.65 0.33 1.17 0.39 1.17 0.39 1.65 0.74 1.65 0.74 1.17 0.8 1.17 0.8 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.565 0.705 1.36 0.705 1.36 0.74 1.24 0.74 1.24 0.625 1.46 0.625 1.46 0.485 1.565 0.485 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.82051275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.865 0.71 0.74 0.71 0.74 0.73 0.66 0.73 0.66 0.67 0.26 0.67 0.26 0.59 0.865 0.59 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.77 0.56 0.9 ;
    END
  END A1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6393 LAYER Metal1 ;
    ANTENNADIFFAREA 1.06325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 1.02 1.205 1.02 1.205 0.9 1.08 0.9 1.08 0.73 1.06 0.73 1.06 0.49 0.575 0.49 0.575 0.47 0.505 0.47 0.505 0.41 0.625 0.41 0.625 0.43 1.08 0.43 1.08 0.37 1.14 0.37 1.14 0.84 1.265 0.84 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      POLYGON 1.47 1.29 0.945 1.29 0.945 1.06 0.595 1.06 0.595 1.29 0.535 1.29 0.535 1.06 0.185 1.06 0.185 1.29 0.125 1.29 0.125 1 1.005 1 1.005 1.23 1.41 1.23 1.41 0.9 1.47 0.9 ;
  END
END AOI21X2

MACRO AOI21X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21X4 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1892 LAYER Metal1 ;
    ANTENNADIFFAREA 1.9498 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.53 1.075 2.47 1.075 2.47 1.015 2.165 1.015 2.165 1.075 2.06 1.075 2.06 0.895 1.89 0.895 1.89 0.525 0.855 0.525 0.855 0.505 0.785 0.505 0.785 0.445 0.905 0.445 0.905 0.465 1.405 0.465 1.405 0.445 1.525 0.445 1.525 0.465 1.95 0.465 1.95 0.405 2.01 0.405 2.01 0.465 2.345 0.465 2.345 0.445 2.465 0.445 2.465 0.505 2.395 0.505 2.395 0.525 1.95 0.525 1.95 0.815 2.165 0.815 2.165 0.955 2.53 0.955 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.0897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 0.815 1.45 0.895 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.75641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 0.92 1.66 0.92 1.66 0.715 0.54 0.715 0.54 0.655 1.74 0.655 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.54 0.715 2.05 0.715 2.05 0.635 2.235 0.635 2.235 0.625 2.365 0.625 2.365 0.635 2.54 0.635 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.77 0 1.77 0 1.65 0.41 1.65 0.41 1.225 0.47 1.225 0.47 1.65 0.82 1.65 0.82 1.225 0.88 1.225 0.88 1.65 1.23 1.65 1.23 1.225 1.29 1.225 1.29 1.65 1.64 1.65 1.64 1.225 1.7 1.225 1.7 1.65 3 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 0.06 2.64 0.06 2.64 0.395 2.58 0.395 2.58 0.06 2.185 0.06 2.185 0.305 2.245 0.305 2.245 0.365 2.125 0.365 2.125 0.06 1.775 0.06 1.775 0.305 1.835 0.305 1.835 0.365 1.715 0.365 1.715 0.06 1.155 0.06 1.155 0.305 1.215 0.305 1.215 0.365 1.095 0.365 1.095 0.06 0.565 0.06 0.565 0.395 0.505 0.395 0.505 0.06 0 0.06 0 -0.06 3 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.735 1.345 1.845 1.345 1.845 1.08 1.495 1.08 1.495 1.345 1.435 1.345 1.435 1.08 1.085 1.08 1.085 1.345 1.025 1.345 1.025 1.08 0.675 1.08 0.675 1.345 0.615 1.345 0.615 1.08 0.265 1.08 0.265 1.345 0.205 1.345 0.205 1.02 1.905 1.02 1.905 1.285 2.265 1.285 2.265 1.115 2.325 1.115 2.325 1.285 2.675 1.285 2.675 0.955 2.735 0.955 ;
  END
END AOI21X4

MACRO AOI21XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21XL 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.425 LAYER Metal1 ;
    ANTENNADIFFAREA 0.490725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 0.73 0.92 0.73 0.92 1.295 0.9 1.295 0.9 1.355 0.84 1.355 0.84 1.235 0.86 1.235 0.86 0.63 0.64 0.63 0.64 0.405 0.7 0.405 0.7 0.57 0.92 0.57 0.92 0.6 0.94 0.6 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.36 0.69 0.14 0.69 0.14 0.88 0.06 0.88 0.06 0.6 0.14 0.6 0.14 0.61 0.36 0.61 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.22 0.54 0.72 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.73 0.74 1.23 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.4 1.65 0.4 1.51 0.46 1.51 0.46 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.875 0.06 0.875 0.41 0.935 0.41 0.935 0.47 0.815 0.47 0.815 0.06 0.305 0.06 0.305 0.5 0.245 0.5 0.245 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.695 1.45 0.615 1.45 0.615 1.41 0.135 1.41 0.135 1.33 0.695 1.33 ;
  END
END AOI21XL

MACRO AOI221X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.64235 LAYER Metal1 ;
    ANTENNADIFFAREA 1.02855 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 1.125 1.315 1.125 1.315 1.3 1.255 1.3 1.255 0.46 0.61 0.46 0.61 0.4 1.235 0.4 1.235 0.22 1.315 0.22 1.315 0.955 1.34 0.955 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.4102565 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.58 0.75 0.92 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.4102565 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.58 0.95 0.92 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.25641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.34 0.575 0.315 0.575 0.315 0.66 0.28 0.66 0.28 0.665 0.185 0.665 0.185 0.53 0.26 0.53 0.26 0.405 0.34 0.405 ;
    END
  END A0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.12820525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 0.58 1.19 0.73 ;
    END
  END C0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.076923 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 0.745 0.385 0.745 0.385 0.62 0.43 0.62 0.43 0.6 0.54 0.6 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.92 0.13 0.92 0.13 1.65 0.51 1.65 0.51 1.385 0.57 1.385 0.57 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 0.99 0.06 0.99 0.26 1.05 0.26 1.05 0.32 0.93 0.32 0.93 0.06 0.165 0.06 0.165 0.47 0.105 0.47 0.105 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.11 1.3 0.64 1.3 0.64 1.18 0.7 1.18 0.7 1.24 1.05 1.24 1.05 0.98 1.11 0.98 ;
      POLYGON 0.935 1.11 0.335 1.11 0.335 1.185 0.275 1.185 0.275 1.05 0.935 1.05 ;
  END
END AOI221X1

MACRO AOI221X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X2 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2359 LAYER Metal1 ;
    ANTENNADIFFAREA 1.7726 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.28 1.135 2.22 1.135 2.22 1.055 1.08 1.055 1.08 0.92 1.06 0.92 1.06 0.79 1.08 0.79 1.08 0.51 0.605 0.51 0.605 0.45 2.17 0.45 2.17 0.51 1.14 0.51 1.14 0.995 2.28 0.995 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 0.815 1.935 0.895 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.765 0.74 1.065 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.25641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.96 0.69 0.365 0.69 0.365 0.715 0.235 0.715 0.235 0.625 0.285 0.625 0.285 0.61 0.96 0.61 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.025641 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.935 0.715 1.24 0.715 1.24 0.635 1.635 0.635 1.635 0.625 1.765 0.625 1.765 0.635 1.935 0.635 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.065 0.815 2.565 0.895 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 1.77 0 1.77 0 1.65 0.125 1.65 0.125 1.015 0.185 1.015 0.185 1.65 0.505 1.65 0.505 1.315 0.625 1.315 0.625 1.375 0.565 1.375 0.565 1.65 0.915 1.65 0.915 1.315 1.035 1.315 1.035 1.375 0.975 1.375 0.975 1.65 2.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 0.06 2.345 0.06 2.345 0.41 2.285 0.41 2.285 0.06 1.875 0.06 1.875 0.29 1.935 0.29 1.935 0.35 1.815 0.35 1.815 0.06 1.005 0.06 1.005 0.29 1.065 0.29 1.065 0.35 0.945 0.35 0.945 0.06 0.385 0.06 0.385 0.41 0.325 0.41 0.325 0.06 0 0.06 0 -0.06 2.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.485 1.435 1.24 1.435 1.24 1.375 1.165 1.375 1.165 1.315 1.3 1.315 1.3 1.375 1.575 1.375 1.575 1.315 1.695 1.315 1.695 1.375 2.015 1.375 2.015 1.285 2.075 1.285 2.075 1.375 2.425 1.375 2.425 1.015 2.485 1.015 ;
      POLYGON 1.87 1.275 1.81 1.275 1.81 1.215 1.46 1.215 1.46 1.275 1.4 1.275 1.4 1.215 0.8 1.215 0.8 1.275 0.74 1.275 0.74 1.215 0.39 1.215 0.39 1.405 0.33 1.405 0.33 1.015 0.39 1.015 0.39 1.155 1.87 1.155 ;
  END
END AOI221X2

MACRO AOI221X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221X4 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2951 LAYER Metal1 ;
    ANTENNADIFFAREA 3.249 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.305 1.135 4.245 1.135 4.245 1.055 3.895 1.055 3.895 1.135 3.835 1.135 3.835 1.055 1.905 1.055 1.905 0.705 1.835 0.705 1.835 0.625 1.905 0.625 1.905 0.525 0.83 0.525 0.83 0.505 0.76 0.505 0.76 0.445 0.88 0.445 0.88 0.465 1.38 0.465 1.38 0.445 1.5 0.445 1.5 0.465 2.37 0.465 2.37 0.445 2.49 0.445 2.49 0.465 3.135 0.465 3.135 0.445 3.255 0.445 3.255 0.465 3.675 0.465 3.675 0.445 3.795 0.445 3.795 0.465 4.115 0.465 4.115 0.445 4.235 0.445 4.235 0.505 4.165 0.505 4.165 0.525 1.965 0.525 1.965 0.995 4.305 0.995 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.102564 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.685 0.815 1.425 0.895 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.5 0.815 3.18 0.895 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.0641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.735 0.705 0.23 0.705 0.23 0.645 0.235 0.645 0.235 0.625 0.365 0.625 0.365 0.645 1.735 0.645 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.551282 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.565 0.895 3.425 0.895 3.425 0.715 2.09 0.715 2.09 0.655 3.545 0.655 3.545 0.715 3.485 0.715 3.485 0.815 3.565 0.815 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.6153845 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.195 0.71 3.965 0.71 3.965 0.895 3.835 0.895 3.835 0.625 3.965 0.625 3.965 0.63 4.195 0.63 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.77 0 1.77 0 1.65 0.13 1.65 0.13 1.015 0.19 1.015 0.19 1.65 0.51 1.65 0.51 1.315 0.63 1.315 0.63 1.375 0.57 1.375 0.57 1.65 0.92 1.65 0.92 1.315 1.04 1.315 1.04 1.375 0.98 1.375 0.98 1.65 1.33 1.65 1.33 1.315 1.45 1.315 1.45 1.375 1.39 1.375 1.39 1.65 1.74 1.65 1.74 1.315 1.86 1.315 1.86 1.375 1.8 1.375 1.8 1.65 4.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 0.06 4.41 0.06 4.41 0.395 4.35 0.395 4.35 0.06 3.955 0.06 3.955 0.305 4.015 0.305 4.015 0.365 3.895 0.365 3.895 0.06 3.515 0.06 3.515 0.305 3.575 0.305 3.575 0.365 3.455 0.365 3.455 0.06 2.84 0.06 2.84 0.305 2.9 0.305 2.9 0.365 2.78 0.365 2.78 0.06 1.75 0.06 1.75 0.305 1.81 0.305 1.81 0.365 1.69 0.365 1.69 0.06 1.13 0.06 1.13 0.305 1.19 0.305 1.19 0.365 1.07 0.365 1.07 0.06 0.54 0.06 0.54 0.395 0.48 0.395 0.48 0.06 0 0.06 0 -0.06 4.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.51 1.435 2.02 1.435 2.02 1.375 1.96 1.375 1.96 1.315 2.08 1.315 2.08 1.375 2.37 1.375 2.37 1.315 2.49 1.315 2.49 1.375 2.78 1.375 2.78 1.315 2.9 1.315 2.9 1.375 3.19 1.375 3.19 1.315 3.31 1.315 3.31 1.375 3.63 1.375 3.63 1.285 3.69 1.285 3.69 1.375 4.04 1.375 4.04 1.155 4.1 1.155 4.1 1.375 4.45 1.375 4.45 1.015 4.51 1.015 ;
      POLYGON 3.485 1.275 3.425 1.275 3.425 1.215 3.075 1.215 3.075 1.275 3.015 1.275 3.015 1.215 2.665 1.215 2.665 1.275 2.605 1.275 2.605 1.215 2.255 1.215 2.255 1.275 2.195 1.275 2.195 1.215 1.625 1.215 1.625 1.405 1.565 1.405 1.565 1.215 1.215 1.215 1.215 1.405 1.155 1.405 1.155 1.215 0.805 1.215 0.805 1.405 0.745 1.405 0.745 1.075 0.395 1.075 0.395 1.405 0.335 1.405 0.335 1.015 0.805 1.015 0.805 1.155 1.155 1.155 1.155 1.015 1.215 1.015 1.215 1.155 1.565 1.155 1.565 1.015 1.625 1.015 1.625 1.155 3.485 1.155 ;
  END
END AOI221X4

MACRO AOI221XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221XL 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8334 LAYER Metal1 ;
    ANTENNADIFFAREA 0.994025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 0.92 1.88 0.92 1.88 1.21 1.82 1.21 1.82 0.7 0.965 0.7 0.965 0.475 1.025 0.475 1.025 0.64 1.715 0.64 1.715 0.475 1.775 0.475 1.775 0.64 1.88 0.64 1.88 0.79 1.94 0.79 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.13 0.955 0.69 0.955 0.69 0.815 0.965 0.815 0.965 0.875 1.13 0.875 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 0.895 1.325 0.895 1.325 1.085 1.245 1.085 1.245 0.895 1.23 0.895 1.23 0.815 1.54 0.815 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.835 0.395 1.085 ;
    END
  END A0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.72 1.085 1.425 1.085 1.425 1.005 1.64 1.005 1.64 0.8 1.72 0.8 ;
    END
  END C0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.9444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.59 0.735 0.47 0.735 0.47 0.325 0.435 0.325 0.435 0.245 0.565 0.245 0.565 0.655 0.59 0.655 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.205 1.65 0.205 1.51 0.265 1.51 0.265 1.65 0.605 1.65 0.605 1.395 0.665 1.395 0.665 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.34 0.06 1.34 0.48 1.4 0.48 1.4 0.54 1.28 0.54 1.28 0.06 0.325 0.06 0.325 0.57 0.265 0.57 0.265 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.445 1.485 0.905 1.485 0.905 1.295 0.865 1.295 0.865 1.215 0.985 1.215 0.985 1.405 1.365 1.405 1.365 1.185 1.445 1.185 ;
      POLYGON 1.23 1.305 1.17 1.305 1.17 1.245 1.085 1.245 1.085 1.115 0.765 1.115 0.765 1.245 0.43 1.245 0.43 1.305 0.37 1.305 0.37 1.185 0.705 1.185 0.705 1.055 1.145 1.055 1.145 1.185 1.23 1.185 ;
  END
END AOI221XL

MACRO AOI222X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X1 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7883 LAYER Metal1 ;
    ANTENNADIFFAREA 1.1808 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 1.26 1.435 1.26 1.435 1.32 1.375 1.32 1.375 1.2 1.66 1.2 1.66 0.52 0.76 0.52 0.76 0.38 0.82 0.38 0.82 0.46 1.45 0.46 1.45 0.41 1.72 0.41 1.72 0.98 1.74 0.98 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 1.1 0.68 1.1 0.68 0.92 0.66 0.92 0.66 0.62 0.76 0.62 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.62 1.54 1.1 ;
    END
  END C1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.49 0.34 0.99 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.095 1.1 0.88 1.1 0.88 0.92 0.86 0.92 0.86 0.755 0.94 0.755 0.94 0.86 1.095 0.86 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.92 1.275 0.92 1.275 1.225 1.195 1.225 1.195 0.79 1.34 0.79 ;
    END
  END C0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.22 0.545 0.715 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.15 1.65 0.15 1.09 0.21 1.09 0.21 1.65 0.56 1.65 0.56 1.36 0.62 1.36 0.62 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.14 0.06 1.14 0.36 1.08 0.36 1.08 0.06 0.31 0.06 0.31 0.36 0.25 0.36 0.25 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.64 1.48 0.76 1.48 0.76 1.36 0.82 1.36 0.82 1.42 1.17 1.42 1.17 1.325 1.23 1.325 1.23 1.42 1.58 1.42 1.58 1.36 1.64 1.36 ;
      POLYGON 1.025 1.32 0.965 1.32 0.965 1.26 0.415 1.26 0.415 1.48 0.355 1.48 0.355 1.2 1.025 1.2 ;
  END
END AOI222X1

MACRO AOI222X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X2 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4936 LAYER Metal1 ;
    ANTENNADIFFAREA 2.1605 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.91 1.135 2.85 1.135 2.85 1.08 2.5 1.08 2.5 1.155 2.44 1.155 2.44 1.065 1.28 1.065 1.28 0.92 1.26 0.92 1.26 0.79 1.28 0.79 1.28 0.51 0.705 0.51 0.705 0.45 2.675 0.45 2.675 0.51 1.34 0.51 1.34 1.005 2.5 1.005 2.5 1.02 2.85 1.02 2.85 1.015 2.91 1.015 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.635 0.815 2.135 0.895 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.5641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.79 0.835 0.92 ;
    END
  END A1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.6153845 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.74 0.895 2.725 0.895 2.725 0.92 2.555 0.92 2.555 0.79 2.725 0.79 2.725 0.815 2.74 0.815 ;
    END
  END C1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.025641 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.06 0.715 0.865 0.715 0.865 0.69 0.56 0.69 0.56 0.74 0.235 0.74 0.235 0.625 0.505 0.625 0.505 0.61 0.95 0.61 0.95 0.635 1.06 0.635 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.69230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.135 0.715 1.505 0.715 1.505 0.635 1.835 0.635 1.835 0.625 1.965 0.625 1.965 0.635 2.135 0.635 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.74358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.015 0.74 2.84 0.74 2.84 0.685 2.4 0.685 2.4 0.715 2.235 0.715 2.235 0.625 2.9 0.625 2.9 0.68 3.015 0.68 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 1.77 0 1.77 0 1.65 0.225 1.65 0.225 1.015 0.285 1.015 0.285 1.65 0.605 1.65 0.605 1.315 0.725 1.315 0.725 1.375 0.665 1.375 0.665 1.65 1.015 1.65 1.015 1.315 1.135 1.315 1.135 1.375 1.075 1.375 1.075 1.65 3.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 0.06 2.955 0.06 2.955 0.435 2.895 0.435 2.895 0.06 2.18 0.06 2.18 0.29 2.24 0.29 2.24 0.35 2.12 0.35 2.12 0.06 1.105 0.06 1.105 0.29 1.165 0.29 1.165 0.35 1.045 0.35 1.045 0.06 0.485 0.06 0.485 0.435 0.425 0.435 0.425 0.06 0 0.06 0 -0.06 3.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.115 1.435 1.435 1.435 1.435 1.375 1.375 1.375 1.375 1.315 1.495 1.315 1.495 1.375 1.795 1.375 1.795 1.315 1.915 1.315 1.915 1.375 2.235 1.375 2.235 1.285 2.295 1.285 2.295 1.375 2.615 1.375 2.615 1.315 2.735 1.315 2.735 1.375 3.055 1.375 3.055 1.015 3.115 1.015 ;
      POLYGON 2.09 1.275 2.03 1.275 2.03 1.215 1.67 1.215 1.67 1.275 1.61 1.275 1.61 1.215 0.9 1.215 0.9 1.405 0.84 1.405 0.84 1.08 0.49 1.08 0.49 1.405 0.43 1.405 0.43 1.015 0.49 1.015 0.49 1.02 0.84 1.02 0.84 1.015 0.9 1.015 0.9 1.155 2.09 1.155 ;
  END
END AOI222X2

MACRO AOI222X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222X4 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6881 LAYER Metal1 ;
    ANTENNADIFFAREA 3.8452 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.145 1.135 5.085 1.135 5.085 1.055 4.735 1.055 4.735 1.135 4.675 1.135 4.675 1.055 4.325 1.055 4.325 1.135 4.265 1.135 4.265 1.055 3.915 1.055 3.915 1.135 3.855 1.135 3.855 1.055 1.905 1.055 1.905 0.895 1.835 0.895 1.835 0.815 1.905 0.815 1.905 0.555 0.83 0.555 0.83 0.535 0.76 0.535 0.76 0.475 0.88 0.475 0.88 0.495 1.38 0.495 1.38 0.475 1.5 0.475 1.5 0.495 2.345 0.495 2.345 0.475 2.465 0.475 2.465 0.495 3.21 0.495 3.21 0.475 3.33 0.475 3.33 0.495 3.98 0.495 3.98 0.475 4.1 0.475 4.1 0.495 4.51 0.495 4.51 0.475 4.72 0.475 4.72 0.535 4.56 0.535 4.56 0.555 1.965 0.555 1.965 0.995 5.145 0.995 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.0897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.465 0.815 3.2 0.895 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.815 1.425 0.895 ;
    END
  END A1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.102564 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.055 0.815 4.795 0.895 ;
    END
  END C1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.64102575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.61 0.715 2.295 0.715 2.295 0.815 2.365 0.815 2.365 0.895 2.235 0.895 2.235 0.715 2.11 0.715 2.11 0.655 3.61 0.655 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.83333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.15 0.715 3.745 0.715 3.745 0.655 4.835 0.655 4.835 0.625 4.965 0.625 4.965 0.655 5.15 0.655 ;
    END
  END C0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.602564 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.735 0.715 0.42 0.715 0.42 0.655 0.435 0.655 0.435 0.625 0.565 0.625 0.565 0.655 1.735 0.655 ;
    END
  END A0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 0 1.77 0 1.65 0.135 1.65 0.135 1.015 0.195 1.015 0.195 1.65 0.515 1.65 0.515 1.315 0.635 1.315 0.635 1.375 0.575 1.375 0.575 1.65 0.925 1.65 0.925 1.315 1.045 1.315 1.045 1.375 0.985 1.375 0.985 1.65 1.335 1.65 1.335 1.315 1.455 1.315 1.455 1.375 1.395 1.375 1.395 1.65 1.745 1.65 1.745 1.315 1.865 1.315 1.865 1.375 1.805 1.375 1.805 1.65 5.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5 0.06 5 0.425 4.94 0.425 4.94 0.06 4.35 0.06 4.35 0.335 4.41 0.335 4.41 0.395 4.29 0.395 4.29 0.06 3.68 0.06 3.68 0.335 3.74 0.335 3.74 0.395 3.62 0.395 3.62 0.06 2.715 0.06 2.715 0.335 2.775 0.335 2.775 0.395 2.655 0.395 2.655 0.06 1.75 0.06 1.75 0.335 1.81 0.335 1.81 0.395 1.69 0.395 1.69 0.06 1.13 0.06 1.13 0.335 1.19 0.335 1.19 0.395 1.07 0.395 1.07 0.06 0.54 0.06 0.54 0.425 0.48 0.425 0.48 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.35 1.435 2.04 1.435 2.04 1.375 1.98 1.375 1.98 1.315 2.1 1.315 2.1 1.375 2.39 1.375 2.39 1.315 2.51 1.315 2.51 1.375 2.8 1.375 2.8 1.315 2.92 1.315 2.92 1.375 3.21 1.375 3.21 1.315 3.33 1.315 3.33 1.375 3.65 1.375 3.65 1.285 3.71 1.285 3.71 1.375 4.06 1.375 4.06 1.285 4.12 1.285 4.12 1.375 4.47 1.375 4.47 1.285 4.53 1.285 4.53 1.375 4.88 1.375 4.88 1.285 4.94 1.285 4.94 1.375 5.29 1.375 5.29 1.015 5.35 1.015 ;
      POLYGON 3.505 1.275 3.445 1.275 3.445 1.215 3.095 1.215 3.095 1.275 3.035 1.275 3.035 1.215 2.685 1.215 2.685 1.275 2.625 1.275 2.625 1.215 2.275 1.215 2.275 1.275 2.215 1.275 2.215 1.215 1.63 1.215 1.63 1.405 1.57 1.405 1.57 1.215 1.22 1.215 1.22 1.405 1.16 1.405 1.16 1.215 0.81 1.215 0.81 1.405 0.75 1.405 0.75 1.215 0.4 1.215 0.4 1.405 0.34 1.405 0.34 1.015 0.4 1.015 0.4 1.155 0.75 1.155 0.75 1.015 0.81 1.015 0.81 1.155 1.16 1.155 1.16 1.015 1.22 1.015 1.22 1.155 1.57 1.155 1.57 1.015 1.63 1.015 1.63 1.155 3.505 1.155 ;
  END
END AOI222X4

MACRO AOI222XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222XL 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8243 LAYER Metal1 ;
    ANTENNADIFFAREA 1.0364 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 0.54 1.92 0.54 1.92 1.07 1.645 1.07 1.645 1.195 1.585 1.195 1.585 1.01 1.86 1.01 1.86 0.33 0.9 0.33 0.9 0.36 0.84 0.36 0.84 0.24 0.9 0.24 0.9 0.27 1.92 0.27 1.92 0.41 1.94 0.41 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.095 0.895 0.835 0.895 0.835 0.575 1.025 0.575 1.025 0.815 1.095 0.815 ;
    END
  END B1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.76 0.91 1.62 0.91 1.62 0.83 1.66 0.83 1.66 0.47 1.74 0.47 1.74 0.83 1.76 0.83 ;
    END
  END C1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.335 0.895 0.035 0.895 0.035 0.815 0.215 0.815 0.215 0.615 0.335 0.615 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 1.035 1.26 1.035 1.26 0.825 1.195 0.825 1.195 0.745 1.26 0.745 1.26 0.6 1.34 0.6 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 0.73 1.52 0.73 1.52 0.91 1.44 0.91 1.44 0.43 1.54 0.43 ;
    END
  END C0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.58 0.895 0.435 0.895 0.435 0.46 0.555 0.46 0.555 0.815 0.58 0.815 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.145 1.65 0.145 1.51 0.205 1.51 0.205 1.65 0.57 1.65 0.57 1.51 0.63 1.51 0.63 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.41 0.06 1.41 0.17 1.29 0.17 1.29 0.06 0.24 0.06 0.24 0.36 0.18 0.36 0.18 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.85 1.29 1.805 1.29 1.805 1.355 0.92 1.355 0.92 1.26 0.86 1.26 0.86 1.2 0.98 1.2 0.98 1.295 1.3 1.295 1.3 1.17 1.36 1.17 1.36 1.295 1.745 1.295 1.745 1.23 1.79 1.23 1.79 1.17 1.85 1.17 ;
      POLYGON 1.16 1.195 1.08 1.195 1.08 1.1 0.415 1.1 0.415 1.14 0.335 1.14 0.335 1.02 1.16 1.02 ;
  END
END AOI222XL

MACRO AOI22X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4692 LAYER Metal1 ;
    ANTENNADIFFAREA 0.7856 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.755 1.325 0.695 1.325 0.695 1.085 0.455 1.085 0.455 0.525 0.485 0.525 0.485 0.23 0.545 0.23 0.545 0.595 0.515 0.595 0.515 1.005 0.755 1.005 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.4358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.55 0.18 0.765 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.897436 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.965 0.735 0.805 0.735 0.805 0.725 0.77 0.725 0.77 0.55 0.965 0.55 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.051282 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 0.93 0.59 0.93 0.59 0.685 0.65 0.685 0.65 0.795 0.74 0.795 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.79487175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.395 0.365 0.66 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.245 1.65 0.245 1.37 0.365 1.37 0.365 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.905 0.06 0.905 0.49 0.845 0.49 0.845 0.06 0.13 0.06 0.13 0.49 0.07 0.49 0.07 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.96 1.46 0.48 1.46 0.48 1.27 0.13 1.27 0.13 1.46 0.07 1.46 0.07 1.21 0.54 1.21 0.54 1.4 0.9 1.4 0.9 1.07 0.96 1.07 ;
  END
END AOI22X1

MACRO AOI22X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X2 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8496 LAYER Metal1 ;
    ANTENNADIFFAREA 1.51965 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.9 1.165 1.43 1.165 1.43 0.895 1.035 0.895 1.035 0.815 1.165 0.815 1.165 0.475 0.71 0.475 0.71 0.415 1.685 0.415 1.685 0.475 1.225 0.475 1.225 0.835 1.49 0.835 1.49 1.105 1.84 1.105 1.84 0.995 1.9 0.995 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.71794875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.655 0.715 0.745 0.96 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.897436 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.74 1.74 1.03 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.30769225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.165 0.895 1.84 0.895 1.84 0.64 1.56 0.64 1.56 0.715 1.325 0.715 1.325 0.655 1.5 0.655 1.5 0.58 1.96 0.58 1.96 0.815 2.165 0.815 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.065 0.715 0.84 0.715 0.84 0.655 0.56 0.655 0.56 0.705 0.235 0.705 0.235 0.625 0.48 0.625 0.48 0.575 0.92 0.575 0.92 0.635 1.065 0.635 ;
    END
  END A0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.345 1.65 0.345 1.195 0.405 1.195 0.405 1.65 0.725 1.65 0.725 1.225 0.845 1.225 0.845 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 2.005 0.06 2.005 0.435 1.945 0.435 1.945 0.06 1.11 0.06 1.11 0.255 1.17 0.255 1.17 0.315 1.05 0.315 1.05 0.06 0.49 0.06 0.49 0.435 0.43 0.435 0.43 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.105 1.285 1.05 1.285 1.05 1.08 0.61 1.08 0.61 1.315 0.55 1.315 0.55 1.08 0.2 1.08 0.2 1.315 0.14 1.315 0.14 0.925 0.2 0.925 0.2 1.02 1.05 1.02 1.05 0.995 1.11 0.995 1.11 1.225 2.045 1.225 2.045 0.995 2.105 0.995 ;
  END
END AOI22X2

MACRO AOI22X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22X4 0 0 ;
  SIZE 3.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3824 LAYER Metal1 ;
    ANTENNADIFFAREA 2.45 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.25 1.115 3.19 1.115 3.19 1.055 2.84 1.055 2.84 1.115 2.78 1.115 2.78 1.055 2.43 1.055 2.43 1.115 2.37 1.115 2.37 1.055 2.02 1.055 2.02 1.115 1.96 1.115 1.96 0.895 1.74 0.895 1.74 0.525 0.765 0.525 0.765 0.505 0.695 0.505 0.695 0.445 0.815 0.445 0.815 0.465 1.315 0.465 1.315 0.445 1.435 0.445 1.435 0.465 2.135 0.465 2.135 0.445 2.255 0.445 2.255 0.465 2.665 0.465 2.665 0.445 2.875 0.445 2.875 0.505 2.715 0.505 2.715 0.525 1.8 0.525 1.8 0.815 1.965 0.815 1.965 0.835 2.02 0.835 2.02 0.995 3.25 0.995 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.0897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.21 0.815 2.945 0.895 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.0897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.625 0.815 1.36 0.895 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.4102565 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.64 0.745 1.54 0.745 1.54 0.92 1.46 0.92 1.46 0.715 0.215 0.715 0.215 0.655 1.58 0.655 1.58 0.625 1.64 0.625 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.9358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.355 0.705 1.9 0.705 1.9 0.645 2.035 0.645 2.035 0.625 2.165 0.625 2.165 0.645 3.355 0.645 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 1.77 0 1.77 0 1.65 0.32 1.65 0.32 1.225 0.38 1.225 0.38 1.65 0.73 1.65 0.73 1.225 0.79 1.225 0.79 1.65 1.14 1.65 1.14 1.225 1.2 1.225 1.2 1.65 1.55 1.65 1.55 1.225 1.61 1.225 1.61 1.65 3.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 0.06 3.155 0.06 3.155 0.395 3.095 0.395 3.095 0.06 2.505 0.06 2.505 0.305 2.565 0.305 2.565 0.365 2.445 0.365 2.445 0.06 1.785 0.06 1.785 0.305 1.845 0.305 1.845 0.365 1.725 0.365 1.725 0.06 1.065 0.06 1.065 0.305 1.125 0.305 1.125 0.365 1.005 0.365 1.005 0.06 0.475 0.06 0.475 0.395 0.415 0.395 0.415 0.06 0 0.06 0 -0.06 3.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.455 1.345 1.755 1.345 1.755 1.08 1.405 1.08 1.405 1.345 1.345 1.345 1.345 1.08 0.995 1.08 0.995 1.345 0.935 1.345 0.935 1.08 0.585 1.08 0.585 1.345 0.525 1.345 0.525 1.08 0.175 1.08 0.175 1.345 0.115 1.345 0.115 1.02 1.815 1.02 1.815 1.285 2.165 1.285 2.165 1.225 2.225 1.225 2.225 1.285 2.575 1.285 2.575 1.225 2.635 1.225 2.635 1.285 2.985 1.285 2.985 1.225 3.045 1.225 3.045 1.285 3.395 1.285 3.395 0.955 3.455 0.955 ;
  END
END AOI22X4

MACRO AOI22XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.521425 LAYER Metal1 ;
    ANTENNADIFFAREA 0.5832 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.805 1.235 0.745 1.235 0.745 1.175 0.7 1.175 0.7 1.11 0.635 1.11 0.635 1.005 0.5 1.005 0.5 0.62 0.52 0.62 0.52 0.255 0.58 0.255 0.58 0.945 0.77 0.945 0.77 1.115 0.805 1.115 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.388889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.18 0.975 0.06 0.975 0.06 0.75 0.155 0.75 0.155 0.785 0.18 0.785 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.388889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.7 0.98 0.925 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.78 0.73 0.68 0.73 0.68 0.515 0.66 0.515 0.66 0.435 0.68 0.435 0.68 0.25 0.76 0.25 0.76 0.53 0.78 0.53 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.9814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.4 0.54 0.365 0.54 0.365 0.73 0.235 0.73 0.235 0.41 0.4 0.41 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.21 0.335 1.21 0.335 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 1.01 0.06 1.01 0.35 0.95 0.35 0.95 0.06 0.13 0.06 0.13 0.35 0.07 0.35 0.07 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.01 1.395 0.48 1.395 0.48 1.15 0.13 1.15 0.13 1.235 0.07 1.235 0.07 1.09 0.54 1.09 0.54 1.335 0.95 1.335 0.95 1.21 1.01 1.21 ;
  END
END AOI22XL

MACRO AOI2BB1X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.477 LAYER Metal1 ;
    ANTENNADIFFAREA 0.642025 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.30769225 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 134.87179475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.49 0.475 0.42 0.475 0.42 0.515 0.235 0.515 0.235 0.755 0.31 0.755 0.31 1.475 0.25 1.475 0.25 0.815 0.175 0.815 0.175 0.435 0.37 0.435 0.37 0.415 0.49 0.415 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.42 0.755 0.56 1.135 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.715 0.74 1.045 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.4814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1 0.58 1.14 0.79 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.56 1.65 0.56 1.21 0.62 1.21 0.62 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 1.105 0.06 1.105 0.48 1.045 0.48 1.045 0.06 0.665 0.06 0.665 0.48 0.605 0.48 0.605 0.06 0.21 0.06 0.21 0.275 0.27 0.275 0.27 0.335 0.15 0.335 0.15 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.005 1.27 0.84 1.27 0.84 0.655 0.295 0.655 0.295 0.595 0.84 0.595 0.84 0.385 0.9 0.385 0.9 1.21 1.005 1.21 ;
  END
END AOI2BB1X1

MACRO AOI2BB1X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8116 LAYER Metal1 ;
    ANTENNADIFFAREA 0.97455 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.87350425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 104.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.9 0.51 0.14 0.51 0.14 1.045 0.695 1.045 0.695 1.43 0.635 1.43 0.635 1.105 0.08 1.105 0.08 0.73 0.06 0.73 0.06 0.6 0.08 0.6 0.08 0.45 0.43 0.45 0.43 0.37 0.49 0.37 0.49 0.45 0.84 0.45 0.84 0.37 0.9 0.37 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.17948725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.96 0.785 0.54 0.785 0.54 0.92 0.46 0.92 0.46 0.785 0.36 0.785 0.36 0.705 0.96 0.705 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.89 1.12 0.89 1.12 0.73 1.06 0.73 1.06 0.45 1.14 0.45 1.14 0.6 1.2 0.6 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.565 1.54 1.065 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.325 1.65 0.325 1.31 0.385 1.31 0.385 1.65 0.945 1.65 0.945 1.15 1.005 1.15 1.005 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.66 0.06 1.66 0.465 1.6 0.465 1.6 0.06 1.105 0.06 1.105 0.35 1.045 0.35 1.045 0.06 0.695 0.06 0.695 0.35 0.635 0.35 0.635 0.06 0.285 0.06 0.285 0.35 0.225 0.35 0.225 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.4 1.225 1.28 1.225 1.28 1.05 0.9 1.05 0.9 0.945 0.67 0.945 0.67 0.885 0.96 0.885 0.96 0.99 1.3 0.99 1.3 0.345 1.36 0.345 1.36 1.165 1.4 1.165 ;
  END
END AOI2BB1X2

MACRO AOI2BB1X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1X4 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.175475 LAYER Metal1 ;
    ANTENNADIFFAREA 1.5887 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.04679475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 75.76923075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.695 0.525 0.235 0.525 0.235 1.195 1.29 1.195 1.29 1.475 1.23 1.475 1.23 1.255 0.67 1.255 0.67 1.475 0.61 1.475 0.61 1.255 0.365 1.255 0.365 1.275 0.235 1.275 0.235 1.255 0.175 1.255 0.175 0.465 0.405 0.465 0.405 0.385 0.465 0.385 0.465 0.465 0.815 0.465 0.815 0.385 0.875 0.385 0.875 0.465 1.225 0.465 1.225 0.385 1.285 0.385 1.285 0.465 1.635 0.465 1.635 0.385 1.695 0.385 ;
    END
  END Y
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.435 1.94 0.935 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.5 2.34 1 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.9871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.755 0.845 0.54 0.845 0.54 0.92 0.46 0.92 0.46 0.845 0.335 0.845 0.335 0.785 1.755 0.785 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 1.77 0 1.77 0 1.65 0.24 1.65 0.24 1.385 0.36 1.385 0.36 1.445 0.3 1.445 0.3 1.65 0.92 1.65 0.92 1.355 0.98 1.355 0.98 1.65 1.74 1.65 1.74 1.195 1.8 1.195 1.8 1.65 2.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 0.06 2.31 0.06 2.31 0.365 2.25 0.365 2.25 0.06 1.93 0.06 1.93 0.335 1.81 0.335 1.81 0.06 1.49 0.06 1.49 0.365 1.43 0.365 1.43 0.06 1.08 0.06 1.08 0.365 1.02 0.365 1.02 0.06 0.67 0.06 0.67 0.365 0.61 0.365 0.61 0.06 0.26 0.06 0.26 0.365 0.2 0.365 0.2 0.06 0 0.06 0 -0.06 2.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.11 1.475 2.05 1.475 2.05 1.095 1.1 1.095 1.1 1.005 0.655 1.005 0.655 0.945 1.16 0.945 1.16 1.035 1.26 1.035 1.26 0.955 1.38 0.955 1.38 1.035 2.045 1.035 2.045 0.385 2.105 0.385 2.105 1.06 2.11 1.06 ;
  END
END AOI2BB1X4

MACRO AOI2BB1XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB1XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4638 LAYER Metal1 ;
    ANTENNADIFFAREA 0.524375 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 28.62962975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 239.35185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.45 0.345 0.375 0.345 0.375 0.51 0.14 0.51 0.14 0.86 0.315 0.86 0.315 1.385 0.255 1.385 0.255 0.92 0.06 0.92 0.06 0.79 0.08 0.79 0.08 0.45 0.315 0.45 0.315 0.285 0.45 0.285 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.55 1.06 0.54 1.06 0.54 1.26 0.46 1.26 0.46 0.98 0.47 0.98 0.47 0.77 0.55 0.77 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 1.26 0.65 1.26 0.65 0.77 0.73 0.77 0.73 0.98 0.74 0.98 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.5555555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 0.84 1.06 0.84 1.06 0.615 0.97 0.615 0.97 0.44 1.03 0.44 1.03 0.54 1.14 0.54 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.565 1.65 0.565 1.36 0.625 1.36 0.625 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 1.06 0.06 1.06 0.35 1 0.35 1 0.06 0.625 0.06 0.625 0.35 0.565 0.35 0.565 0.06 0.215 0.06 0.215 0.35 0.155 0.35 0.155 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.975 1.355 0.84 1.355 0.84 0.67 0.29 0.67 0.29 0.61 0.84 0.61 0.84 0.51 0.795 0.51 0.795 0.255 0.855 0.255 0.855 0.45 0.9 0.45 0.9 1.295 0.975 1.295 ;
  END
END AOI2BB1XL

MACRO AOI2BB2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X1 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 0.73 1.88 0.73 1.88 0.92 1.8 0.92 1.8 0.6 1.86 0.6 1.86 0.48 1.94 0.48 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.45 1.54 0.95 ;
    END
  END B1
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 1.02 0.34 1.02 0.34 1.11 0.26 1.11 0.26 0.94 0.47 0.94 0.47 0.83 0.56 0.83 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 0.73 0.34 0.73 0.34 0.84 0.26 0.84 0.26 0.65 0.46 0.65 0.46 0.54 0.54 0.54 ;
    END
  END A1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8934 LAYER Metal1 ;
    ANTENNADIFFAREA 1.2368 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 15.27179475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 121.25641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.7 1.06 1.64 1.06 1.64 0.35 1.405 0.35 1.405 0.245 1.46 0.245 1.46 0.22 1.54 0.22 1.54 0.29 1.7 0.29 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.335 1.65 0.335 1.21 0.395 1.21 0.395 1.65 1.17 1.65 1.17 1.21 1.23 1.21 1.23 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.86 0.06 1.86 0.38 1.8 0.38 1.8 0.06 1.065 0.06 1.065 0.38 1.005 0.38 1.005 0.06 0.425 0.06 0.425 0.2 0.365 0.2 0.365 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.905 1.33 1.375 1.33 1.375 1.11 1.025 1.11 1.025 1.33 0.965 1.33 0.965 1.05 1.435 1.05 1.435 1.27 1.845 1.27 1.845 1.02 1.905 1.02 ;
      POLYGON 1.36 0.69 1.245 0.69 1.245 0.54 0.845 0.54 0.845 0.44 0.16 0.44 0.16 1.235 0.1 1.235 0.1 0.38 0.905 0.38 0.905 0.48 1.305 0.48 1.305 0.57 1.36 0.57 ;
      POLYGON 1.145 0.7 0.745 0.7 0.745 1.18 0.605 1.18 0.605 1.24 0.545 1.24 0.545 1.12 0.685 1.12 0.685 0.54 0.745 0.54 0.745 0.64 1.145 0.64 ;
  END
END AOI2BB2X1

MACRO AOI2BB2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X2 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3932 LAYER Metal1 ;
    ANTENNADIFFAREA 1.83705 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.90769225 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 90.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.57 1.135 2.51 1.135 2.51 1.055 2.16 1.055 2.16 1.135 2.1 1.135 2.1 1.055 1.88 1.055 1.88 0.92 1.86 0.92 1.86 0.79 1.88 0.79 1.88 0.525 1.61 0.525 1.61 0.505 1.405 0.505 1.405 0.445 1.67 0.445 1.67 0.465 2.275 0.465 2.275 0.445 2.395 0.445 2.395 0.505 2.335 0.505 2.335 0.525 1.94 0.525 1.94 0.995 2.57 0.995 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.075 0.805 2.565 0.895 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.4358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.04 0.625 2.63 0.705 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.6 0.54 1.1 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.46 0.34 0.96 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.77 0 1.77 0 1.65 0.44 1.65 0.44 1.32 0.5 1.32 0.5 1.65 1.23 1.65 1.23 1.285 1.29 1.285 1.29 1.65 1.61 1.65 1.61 1.315 1.73 1.315 1.73 1.375 1.67 1.375 1.67 1.65 3 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 0.06 2.675 0.06 2.675 0.395 2.615 0.395 2.615 0.06 1.83 0.06 1.83 0.305 1.89 0.305 1.89 0.365 1.77 0.365 1.77 0.06 1.185 0.06 1.185 0.395 1.125 0.395 1.125 0.06 0.375 0.06 0.375 0.2 0.315 0.2 0.315 0.06 0 0.06 0 -0.06 3 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.775 1.295 1.855 1.295 1.855 1.275 1.845 1.275 1.845 1.215 1.595 1.215 1.595 1.185 1.495 1.185 1.495 1.405 1.435 1.405 1.435 1.185 1.085 1.185 1.085 1.245 1.025 1.245 1.025 1.125 1.655 1.125 1.655 1.155 1.905 1.155 1.905 1.235 2.305 1.235 2.305 1.175 2.365 1.175 2.365 1.235 2.715 1.235 2.715 1.015 2.775 1.015 ;
      POLYGON 1.76 0.845 0.7 0.845 0.7 1.055 0.64 1.055 0.64 0.54 0.7 0.54 0.7 0.785 1.76 0.785 ;
      POLYGON 1.45 0.685 0.8 0.685 0.8 0.36 0.16 0.36 0.16 1.06 0.295 1.06 0.295 1.12 0.1 1.12 0.1 0.3 0.86 0.3 0.86 0.625 1.45 0.625 ;
  END
END AOI2BB2X2

MACRO AOI2BB2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2X4 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2787 LAYER Metal1 ;
    ANTENNADIFFAREA 3.0036 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.234 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.73803425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 75.84615375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.955 1.115 3.895 1.115 3.895 1.055 3.545 1.055 3.545 1.115 3.485 1.115 3.485 1.055 3.135 1.055 3.135 1.115 3.075 1.115 3.075 1.055 2.765 1.055 2.765 1.115 2.665 1.115 2.665 1.085 2.635 1.085 2.635 0.865 2.475 0.865 2.475 0.525 1.47 0.525 1.47 0.505 1.4 0.505 1.4 0.445 1.52 0.445 1.52 0.465 2.02 0.465 2.02 0.445 2.14 0.445 2.14 0.465 2.65 0.465 2.65 0.445 2.99 0.445 2.99 0.505 2.7 0.505 2.7 0.525 2.535 0.525 2.535 0.805 2.695 0.805 2.695 0.995 3.725 0.995 3.725 0.505 3.66 0.505 3.66 0.445 3.785 0.445 3.785 0.995 3.955 0.995 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.8846155 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.97 0.815 3.625 0.895 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.69230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.06 0.7 3.885 0.7 3.885 0.345 3.56 0.345 3.56 0.705 2.635 0.705 2.635 0.625 2.765 0.625 2.765 0.645 3.5 0.645 3.5 0.285 3.945 0.285 3.945 0.64 4.06 0.64 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.695 0.54 1.195 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.695 0.34 1.195 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.405 1.65 0.405 1.295 0.465 1.295 0.465 1.65 1.025 1.65 1.025 1.125 1.085 1.125 1.085 1.65 1.435 1.65 1.435 1.125 1.495 1.125 1.495 1.65 1.845 1.65 1.845 1.125 1.905 1.125 1.905 1.65 2.225 1.65 2.225 1.255 2.345 1.255 2.345 1.315 2.285 1.315 2.285 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 4.105 0.06 4.105 0.395 4.045 0.395 4.045 0.06 3.34 0.06 3.34 0.395 3.28 0.395 3.28 0.06 2.49 0.06 2.49 0.305 2.55 0.305 2.55 0.365 2.43 0.365 2.43 0.06 1.77 0.06 1.77 0.305 1.83 0.305 1.83 0.365 1.71 0.365 1.71 0.06 1.18 0.06 1.18 0.395 1.12 0.395 1.12 0.06 0.39 0.06 0.39 0.435 0.33 0.435 0.33 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.16 1.345 2.46 1.345 2.46 1.025 2.11 1.025 2.11 1.345 2.05 1.345 2.05 1.025 1.7 1.025 1.7 1.345 1.64 1.345 1.64 1.025 1.29 1.025 1.29 1.345 1.23 1.345 1.23 1.025 0.88 1.025 0.88 1.345 0.82 1.345 0.82 0.965 2.52 0.965 2.52 1.285 2.87 1.285 2.87 1.225 2.93 1.225 2.93 1.285 3.28 1.285 3.28 1.225 3.34 1.225 3.34 1.285 3.69 1.285 3.69 1.225 3.75 1.225 3.75 1.285 4.1 1.285 4.1 0.955 4.16 0.955 ;
      POLYGON 2.375 0.845 0.71 0.845 0.71 1.145 0.64 1.145 0.64 1.025 0.65 1.025 0.65 0.455 0.71 0.455 0.71 0.785 2.375 0.785 ;
      POLYGON 2.065 0.685 0.96 0.685 0.96 0.355 0.55 0.355 0.55 0.595 0.16 0.595 0.16 1.295 0.26 1.295 0.26 1.415 0.2 1.415 0.2 1.355 0.1 1.355 0.1 0.535 0.125 0.535 0.125 0.455 0.185 0.455 0.185 0.535 0.49 0.535 0.49 0.295 1.02 0.295 1.02 0.625 2.065 0.625 ;
  END
END AOI2BB2X4

MACRO AOI2BB2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI2BB2XL 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.17 0.895 1.95 0.895 1.95 0.935 1.87 0.935 1.87 0.655 1.95 0.655 1.95 0.815 2.17 0.815 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.61 0.835 1.53 0.835 1.53 0.705 1.24 0.705 1.24 0.625 1.61 0.625 ;
    END
  END B1
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.565 0.91 0.475 0.91 0.475 0.54 0.435 0.54 0.435 0.46 0.565 0.46 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.64 0.34 1.14 ;
    END
  END A1N
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0424 LAYER Metal1 ;
    ANTENNADIFFAREA 1.050275 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 32.1728395 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 246.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.83 1.095 1.71 1.095 1.71 0.525 1.14 0.525 1.14 0.73 1.06 0.73 1.06 0.6 1.08 0.6 1.08 0.465 1.77 0.465 1.77 1.035 1.83 1.035 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.41 1.65 0.41 1.24 0.47 1.24 0.47 1.65 1.28 1.65 1.28 1.095 1.34 1.095 1.34 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 2.005 0.06 2.005 0.555 1.945 0.555 1.945 0.06 1.235 0.06 1.235 0.17 1.115 0.17 1.115 0.06 0.43 0.06 0.43 0.2 0.37 0.2 0.37 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.05 1.185 1.99 1.185 1.99 1.255 1.515 1.255 1.515 1.09 1.455 1.09 1.455 0.995 1.135 0.995 1.135 1.12 1.075 1.12 1.075 0.935 1.515 0.935 1.515 1.03 1.575 1.03 1.575 1.195 1.93 1.195 1.93 1.125 2.05 1.125 ;
      POLYGON 1.5 0.355 1.395 0.355 1.395 0.36 0.265 0.36 0.265 0.54 0.16 0.54 0.16 1.24 0.265 1.24 0.265 1.36 0.205 1.36 0.205 1.3 0.1 1.3 0.1 0.48 0.205 0.48 0.205 0.3 1.335 0.3 1.335 0.295 1.5 0.295 ;
      POLYGON 0.96 0.755 0.9 0.755 0.9 0.695 0.725 0.695 0.725 1.07 0.68 1.07 0.68 1.32 0.62 1.32 0.62 1.01 0.665 1.01 0.665 0.475 0.785 0.475 0.785 0.535 0.725 0.535 0.725 0.635 0.96 0.635 ;
  END
END AOI2BB2XL

MACRO AOI31X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56875 LAYER Metal1 ;
    ANTENNADIFFAREA 0.75145 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.315 1.05 1.315 1.05 1.48 0.99 1.48 0.99 1.2 1.01 1.2 1.01 0.59 0.73 0.59 0.73 0.23 0.79 0.23 0.79 0.53 1.07 0.53 1.07 1.15 1.14 1.15 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.5641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.55 0.34 0.915 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.17948725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 1.11 0.84 1.11 0.84 0.705 0.92 0.705 0.92 0.98 0.94 0.98 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.4102565 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.705 0.74 1.045 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.5641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.55 1.045 0.47 1.045 0.47 0.895 0.46 0.895 0.46 0.815 0.47 0.815 0.47 0.495 0.55 0.495 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.155 1.65 0.155 1.09 0.215 1.09 0.215 1.65 0.565 1.65 0.565 1.24 0.625 1.24 0.625 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.995 0.06 0.995 0.47 0.935 0.47 0.935 0.06 0.315 0.06 0.315 0.47 0.255 0.47 0.255 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.83 1.48 0.77 1.48 0.77 1.33 0.72 1.33 0.72 1.18 0.42 1.18 0.42 1.48 0.36 1.48 0.36 1.12 0.78 1.12 0.78 1.2 0.83 1.2 ;
  END
END AOI31X1

MACRO AOI31X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7956 LAYER Metal1 ;
    ANTENNADIFFAREA 1.3833 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.565 1.065 1.505 1.065 1.505 1.005 1.48 1.005 1.48 0.73 1.46 0.73 1.46 0.6 1.48 0.6 1.48 0.395 0.7 0.395 0.7 0.335 1.48 0.335 1.48 0.275 1.54 0.275 1.54 0.945 1.565 0.945 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.35897425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.715 0.815 1.055 0.935 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.84615375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.055 0.715 0.54 0.715 0.54 0.92 0.46 0.92 0.46 0.715 0.375 0.715 0.375 0.655 1.055 0.655 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.69230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.73 1.155 0.73 1.155 0.555 0.275 0.555 0.275 0.695 0.215 0.695 0.215 0.495 1.215 0.495 1.215 0.6 1.34 0.6 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.495 1.94 0.995 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.215 0.335 1.215 0.335 1.65 0.685 1.65 0.685 1.215 0.745 1.215 0.745 1.65 1.095 1.65 1.095 1.215 1.155 1.215 1.155 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.745 0.06 1.745 0.395 1.685 0.395 1.685 0.06 1.335 0.06 1.335 0.17 1.215 0.17 1.215 0.06 0.2 0.06 0.2 0.305 0.26 0.305 0.26 0.365 0.14 0.365 0.14 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.77 1.335 1.3 1.335 1.3 1.095 0.95 1.095 0.95 1.335 0.89 1.335 0.89 1.095 0.54 1.095 0.54 1.335 0.48 1.335 0.48 1.08 0.13 1.08 0.13 1.335 0.07 1.335 0.07 0.945 0.13 0.945 0.13 1.02 0.54 1.02 0.54 1.035 1.3 1.035 1.3 0.945 1.36 0.945 1.36 1.275 1.71 1.275 1.71 1.095 1.77 1.095 ;
  END
END AOI31X2

MACRO AOI31X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31X4 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.95145 LAYER Metal1 ;
    ANTENNADIFFAREA 2.7164 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.61 0.675 3.52 0.675 3.52 0.98 3.54 0.98 3.54 1.11 3.47 1.11 3.47 1.115 3.41 1.115 3.41 1.055 3.005 1.055 3.005 1.115 2.945 1.115 2.945 0.995 3.46 0.995 3.46 0.675 1.91 0.675 1.91 0.535 1.97 0.535 1.97 0.615 2.32 0.615 2.32 0.535 2.38 0.535 2.38 0.615 2.73 0.615 2.73 0.535 2.79 0.535 2.79 0.615 3.14 0.615 3.14 0.535 3.2 0.535 3.2 0.615 3.55 0.615 3.55 0.535 3.61 0.535 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.69230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.845 0.895 0.435 0.895 0.435 0.775 0.385 0.775 0.385 0.695 0.515 0.695 0.515 0.815 0.845 0.815 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.69230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.665 0.885 1.365 0.885 1.365 0.895 1.205 0.895 1.205 0.695 1.325 0.695 1.325 0.805 1.665 0.805 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.36 0.855 3.165 0.855 3.165 0.895 3.035 0.895 3.035 0.855 2.9 0.855 2.9 0.775 3.36 0.775 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.035 0.815 2.535 0.895 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 1.77 0 1.77 0 1.65 0.485 1.65 0.485 1.225 0.545 1.225 0.545 1.65 0.895 1.65 0.895 1.225 0.955 1.225 0.955 1.65 1.305 1.65 1.305 1.225 1.365 1.225 1.365 1.65 1.715 1.65 1.715 1.225 1.775 1.225 1.775 1.65 2.125 1.65 2.125 1.225 2.185 1.225 2.185 1.65 2.535 1.65 2.535 1.225 2.595 1.225 2.595 1.65 3.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 0.06 3.405 0.06 3.405 0.515 3.345 0.515 3.345 0.06 2.995 0.06 2.995 0.515 2.935 0.515 2.935 0.06 0.745 0.06 0.745 0.435 0.685 0.435 0.685 0.06 0.335 0.06 0.335 0.435 0.275 0.435 0.275 0.06 0 0.06 0 -0.06 3.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.7 1.345 2.74 1.345 2.74 1.055 2.39 1.055 2.39 1.345 2.33 1.345 2.33 1.055 1.98 1.055 1.98 1.345 1.92 1.345 1.92 1.055 1.57 1.055 1.57 1.345 1.51 1.345 1.51 1.055 1.16 1.055 1.16 1.345 1.1 1.345 1.1 1.055 0.75 1.055 0.75 1.345 0.69 1.345 0.69 1.055 0.34 1.055 0.34 1.345 0.28 1.345 0.28 0.995 2.8 0.995 2.8 1.285 3.15 1.285 3.15 1.225 3.21 1.225 3.21 1.285 3.64 1.285 3.64 0.955 3.7 0.955 ;
      POLYGON 2.585 0.515 2.525 0.515 2.525 0.355 2.175 0.355 2.175 0.515 2.115 0.515 2.115 0.355 1.565 0.355 1.565 0.435 1.505 0.435 1.505 0.355 1.155 0.355 1.155 0.435 1.095 0.435 1.095 0.295 2.585 0.295 ;
      POLYGON 1.77 0.595 0.07 0.595 0.07 0.455 0.13 0.455 0.13 0.535 0.48 0.535 0.48 0.455 0.54 0.455 0.54 0.535 0.89 0.535 0.89 0.455 0.95 0.455 0.95 0.535 1.3 0.535 1.3 0.455 1.36 0.455 1.36 0.535 1.71 0.535 1.71 0.455 1.77 0.455 ;
  END
END AOI31X4

MACRO AOI31XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI31XL 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.60785 LAYER Metal1 ;
    ANTENNADIFFAREA 0.78065 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 0.92 1.325 0.92 1.325 1.21 1.265 1.21 1.265 0.795 0.9 0.795 0.9 0.54 0.96 0.54 0.96 0.735 1.325 0.735 1.325 0.79 1.54 0.79 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.34 1.085 0.26 1.085 0.26 0.895 0.055 0.895 0.055 0.79 0.34 0.79 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.165 1.38 1.085 1.38 1.085 1.085 1.035 1.085 1.035 0.93 1.165 0.93 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.085 0.72 1.085 0.72 0.92 0.66 0.92 0.66 0.645 0.8 0.645 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.545 0.91 0.54 0.91 0.54 0.92 0.46 0.92 0.46 0.79 0.465 0.79 0.465 0.425 0.545 0.425 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.175 1.65 0.175 1.51 0.235 1.51 0.235 1.65 0.645 1.65 0.645 1.51 0.705 1.51 0.705 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.165 0.06 1.165 0.635 1.105 0.635 1.105 0.06 0.265 0.06 0.265 0.635 0.205 0.635 0.205 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.94 1.305 0.86 1.305 0.86 1.265 0.38 1.265 0.38 1.185 0.94 1.185 ;
  END
END AOI31XL

MACRO AOI32X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5484 LAYER Metal1 ;
    ANTENNADIFFAREA 0.9516 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.97 1.315 0.91 1.315 0.91 1.085 0.655 1.085 0.655 0.365 0.715 0.365 0.715 1.005 0.97 1.005 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.87179475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.265 0.54 0.365 0.915 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.5384615 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.815 0.475 0.91 0.92 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.5128205 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.475 0.54 0.555 0.9 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.3846155 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.055 0.675 1.135 0.925 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.076923 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.065 0.67 0.145 1.085 ;
    END
  END A0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.185 0.13 1.185 0.13 1.65 0.48 1.65 0.48 1.345 0.54 1.345 0.54 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 1.15 0.06 1.15 0.61 1.09 0.61 1.09 0.06 0.13 0.06 0.13 0.61 0.07 0.61 0.07 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.175 1.465 0.685 1.465 0.685 1.245 0.335 1.245 0.335 1.465 0.275 1.465 0.275 1.185 0.745 1.185 0.745 1.405 1.115 1.405 1.115 1.075 1.175 1.075 ;
  END
END AOI32X1

MACRO AOI32X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X2 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.969 LAYER Metal1 ;
    ANTENNADIFFAREA 1.87055 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.225 2.14 1.225 2.14 1.165 1.79 1.165 1.79 1.225 1.73 1.225 1.73 1.065 1.565 1.065 1.565 1.085 1.435 1.085 1.435 1.005 1.505 1.005 1.505 0.495 0.815 0.495 0.815 0.435 2.025 0.435 2.025 0.495 1.565 0.495 1.565 1.005 1.79 1.005 1.79 1.105 2.2 1.105 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.025641 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.855 0.995 0.6 0.995 0.6 1.085 0.435 1.085 0.435 1.005 0.52 1.005 0.52 0.915 0.855 0.915 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.025641 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 0.92 1.06 0.92 1.06 0.815 0.52 0.815 0.52 0.755 1.14 0.755 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.89 0.875 2.34 1.005 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.025641 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.82 1.26 0.82 1.26 0.655 0.42 0.655 0.42 0.82 0.36 0.82 0.36 0.595 1.34 0.595 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.84615375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.535 0.8 2.415 0.8 2.415 0.705 1.79 0.705 1.79 0.8 1.665 0.8 1.665 0.625 2.535 0.625 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 1.77 0 1.77 0 1.65 0.39 1.65 0.39 1.345 0.51 1.345 0.51 1.405 0.45 1.405 0.45 1.65 0.8 1.65 0.8 1.345 0.92 1.345 0.92 1.405 0.86 1.405 0.86 1.65 1.21 1.65 1.21 1.345 1.33 1.345 1.33 1.405 1.27 1.405 1.27 1.65 2.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 0.06 2.5 0.06 2.5 0.52 2.44 0.52 2.44 0.06 1.48 0.06 1.48 0.16 1.54 0.16 1.54 0.22 1.42 0.22 1.42 0.06 0.345 0.06 0.345 0.43 0.405 0.43 0.405 0.49 0.285 0.49 0.285 0.06 0 0.06 0 -0.06 2.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.5 1.385 1.445 1.385 1.445 1.245 1.095 1.245 1.095 1.435 1.035 1.435 1.035 1.245 0.685 1.245 0.685 1.305 0.625 1.305 0.625 1.245 0.275 1.245 0.275 1.435 0.215 1.435 0.215 1.045 0.275 1.045 0.275 1.185 1.035 1.185 1.035 1.045 1.095 1.045 1.095 1.185 1.505 1.185 1.505 1.325 1.935 1.325 1.935 1.265 1.995 1.265 1.995 1.325 2.44 1.325 2.44 1.045 2.5 1.045 ;
  END
END AOI32X2

MACRO AOI32X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32X4 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7364 LAYER Metal1 ;
    ANTENNADIFFAREA 3.27375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.16 1.115 4.1 1.115 4.1 1.055 3.75 1.055 3.75 1.115 3.69 1.115 3.69 1.055 3.34 1.055 3.34 1.115 3.28 1.115 3.28 1.055 2.965 1.055 2.965 1.115 2.87 1.115 2.87 0.895 2.64 0.895 2.64 0.395 0.835 0.395 0.835 0.335 3.845 0.335 3.845 0.395 2.7 0.395 2.7 0.815 2.965 0.815 2.965 0.995 4.16 0.995 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.4358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.915 0.985 1.11 0.985 1.11 0.895 0.855 0.895 0.855 0.815 1.165 0.815 1.165 0.835 1.17 0.835 1.17 0.925 1.855 0.925 1.855 0.815 1.915 0.815 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.0897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.12 0.815 3.855 0.895 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.82051275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.32 0.715 1.735 0.715 1.735 0.825 1.27 0.825 1.27 0.715 0.74 0.715 0.74 0.92 0.66 0.92 0.66 0.715 0.535 0.715 0.535 0.655 1.33 0.655 1.33 0.765 1.675 0.765 1.675 0.655 2.32 0.655 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.897436 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.54 0.73 2.46 0.73 2.46 0.715 2.42 0.715 2.42 0.655 2.46 0.655 2.46 0.555 1.55 0.555 1.55 0.665 1.43 0.665 1.43 0.555 0.435 0.555 0.435 0.695 0.375 0.695 0.375 0.495 2.52 0.495 2.52 0.6 2.54 0.6 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.9615385 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.265 0.705 2.8 0.705 2.8 0.625 3.165 0.625 3.165 0.645 4.265 0.645 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.77 0 1.77 0 1.65 0.335 1.65 0.335 1.245 0.395 1.245 0.395 1.65 0.745 1.65 0.745 1.245 0.805 1.245 0.805 1.65 1.175 1.65 1.175 1.245 1.235 1.245 1.235 1.65 1.6 1.65 1.6 1.245 1.66 1.245 1.66 1.65 2.01 1.65 2.01 1.245 2.07 1.245 2.07 1.65 2.42 1.65 2.42 1.245 2.48 1.245 2.48 1.65 4.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 0.06 4.125 0.06 4.125 0.395 4.065 0.395 4.065 0.06 3.505 0.06 3.505 0.17 3.385 0.17 3.385 0.06 2.7 0.06 2.7 0.17 2.58 0.17 2.58 0.06 1.455 0.06 1.455 0.17 1.335 0.17 1.335 0.06 0.36 0.06 0.36 0.305 0.42 0.305 0.42 0.365 0.3 0.365 0.3 0.06 0 0.06 0 -0.06 4.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.365 1.365 2.625 1.365 2.625 1.055 2.275 1.055 2.275 1.365 2.215 1.365 2.215 1.145 1.865 1.145 1.865 1.365 1.805 1.365 1.805 1.145 1.455 1.145 1.455 1.365 1.395 1.365 1.395 1.145 1.01 1.145 1.01 1.365 0.95 1.365 0.95 1.145 0.6 1.145 0.6 1.365 0.54 1.365 0.54 1.08 0.19 1.08 0.19 1.365 0.13 1.365 0.13 0.975 0.19 0.975 0.19 1.02 0.6 1.02 0.6 1.085 0.95 1.085 0.95 0.995 1.01 0.995 1.01 1.085 2.215 1.085 2.215 0.975 2.275 0.975 2.275 0.995 2.685 0.995 2.685 1.305 3.075 1.305 3.075 1.245 3.135 1.245 3.135 1.305 3.485 1.305 3.485 1.245 3.545 1.245 3.545 1.305 3.895 1.305 3.895 1.245 3.955 1.245 3.955 1.305 4.305 1.305 4.305 0.975 4.365 0.975 ;
  END
END AOI32X4

MACRO AOI32XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI32XL 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5352 LAYER Metal1 ;
    ANTENNADIFFAREA 0.8003 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.26 1.245 1.2 1.245 1.2 1.11 0.86 1.11 0.86 0.98 0.88 0.98 0.88 0.425 0.94 0.425 0.94 1.05 1.26 1.05 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 0.89 0.48 0.89 0.48 0.54 0.46 0.54 0.46 0.41 0.54 0.41 0.54 0.48 0.56 0.48 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.23 1.14 0.73 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.745 0.715 0.665 0.715 0.665 0.35 0.66 0.35 0.66 0.22 0.74 0.22 0.74 0.27 0.745 0.27 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.44 1.12 1.36 1.12 1.36 0.92 1.26 0.92 1.26 0.72 1.34 0.72 1.34 0.84 1.44 0.84 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.62 0.34 1.12 ;
    END
  END A0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.19 1.65 0.19 1.51 0.25 1.51 0.25 1.65 0.66 1.65 0.66 1.51 0.72 1.51 0.72 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.365 0.06 1.365 0.52 1.305 0.52 1.305 0.06 0.28 0.06 0.28 0.52 0.22 0.52 0.22 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.465 1.34 1.42 1.34 1.42 1.405 0.825 1.405 0.825 1.28 0.395 1.28 0.395 1.22 0.885 1.22 0.885 1.345 1.36 1.345 1.36 1.28 1.405 1.28 1.405 1.22 1.465 1.22 ;
  END
END AOI32XL

MACRO AOI33X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X1 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7794 LAYER Metal1 ;
    ANTENNADIFFAREA 1.07625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 1.2 1.52 1.2 1.52 1.48 1.46 1.48 1.46 1.18 1.06 1.18 1.06 1.345 1 1.345 1 1.18 0.96 1.18 0.96 1.12 1.46 1.12 1.46 0.61 1.085 0.61 1.085 0.5 0.795 0.5 0.795 0.25 0.855 0.25 0.855 0.44 1.155 0.44 1.155 0.55 1.52 0.55 1.52 1.12 1.54 1.12 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.55 0.34 0.99 ;
    END
  END A0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.645 0.25 0.725 0.75 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.5641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.155 0.87 1.14 0.87 1.14 1.02 1.06 1.02 1.06 0.79 1.075 0.79 1.075 0.67 1.155 0.67 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.82051275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.67 1.34 1.06 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.345 0.54 0.845 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.12820525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 0.94 1.02 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.145 1.65 0.145 1.09 0.205 1.09 0.205 1.65 0.555 1.65 0.555 1.24 0.615 1.24 0.615 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.4 0.06 1.4 0.49 1.28 0.49 1.28 0.06 0.305 0.06 0.305 0.49 0.245 0.49 0.245 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.265 1.48 0.76 1.48 0.76 1.18 0.41 1.18 0.41 1.48 0.35 1.48 0.35 1.09 0.41 1.09 0.41 1.12 0.82 1.12 0.82 1.42 1.205 1.42 1.205 1.24 1.265 1.24 ;
  END
END AOI33X1

MACRO AOI33X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X2 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0953 LAYER Metal1 ;
    ANTENNADIFFAREA 2.1716 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.65 1.165 2.59 1.165 2.59 1.105 2.22 1.105 2.22 1.165 2.16 1.165 2.16 1.105 1.795 1.105 1.795 1.165 1.735 1.165 1.735 1.085 1.435 1.085 1.435 1.005 1.5 1.005 1.5 0.395 0.755 0.395 0.755 0.335 2.195 0.335 2.195 0.395 1.56 0.395 1.56 1.005 1.565 1.005 1.565 1.025 1.795 1.025 1.795 1.045 2.65 1.045 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.16 0.895 0.965 0.895 0.965 0.92 0.685 0.92 0.685 0.815 1.16 0.815 ;
    END
  END A2
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.36 0.895 2.14 0.895 2.14 0.93 1.895 0.93 1.895 0.815 2.36 0.815 ;
    END
  END B2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.54 0.92 2.46 0.92 2.46 0.715 1.84 0.715 1.84 0.655 2.54 0.655 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.897436 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.11 0.715 0.54 0.715 0.54 0.92 0.46 0.92 0.46 0.715 0.42 0.715 0.42 0.655 1.11 0.655 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.64102575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.735 1.26 0.735 1.26 0.555 0.32 0.555 0.32 0.725 0.26 0.725 0.26 0.495 1.32 0.495 1.32 0.6 1.34 0.6 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.7 0.735 2.64 0.735 2.64 0.555 1.74 0.555 1.74 0.735 1.66 0.735 1.66 0.6 1.68 0.6 1.68 0.495 2.7 0.495 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.77 0 1.77 0 1.65 0.29 1.65 0.29 1.345 0.41 1.345 0.41 1.405 0.35 1.405 0.35 1.65 0.7 1.65 0.7 1.345 0.82 1.345 0.82 1.405 0.76 1.405 0.76 1.65 1.11 1.65 1.11 1.345 1.23 1.345 1.23 1.405 1.17 1.405 1.17 1.65 3 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 0.06 2.745 0.06 2.745 0.335 2.805 0.335 2.805 0.395 2.685 0.395 2.685 0.06 1.51 0.06 1.51 0.17 1.39 0.17 1.39 0.06 0.245 0.06 0.245 0.335 0.305 0.335 0.305 0.395 0.185 0.395 0.185 0.06 0 0.06 0 -0.06 3 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.855 1.325 1.39 1.325 1.39 1.245 0.995 1.245 0.995 1.435 0.935 1.435 0.935 1.245 0.585 1.245 0.585 1.435 0.525 1.435 0.525 1.245 0.175 1.245 0.175 1.435 0.115 1.435 0.115 1.045 0.175 1.045 0.175 1.185 0.525 1.185 0.525 1.045 0.585 1.045 0.585 1.185 0.935 1.185 0.935 1.045 0.995 1.045 0.995 1.185 1.45 1.185 1.45 1.265 1.945 1.265 1.945 1.205 2.005 1.205 2.005 1.265 2.365 1.265 2.365 1.205 2.425 1.205 2.425 1.265 2.795 1.265 2.795 1.045 2.855 1.045 ;
  END
END AOI33X2

MACRO AOI33X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33X4 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9833 LAYER Metal1 ;
    ANTENNADIFFAREA 3.91945 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.08 1.205 5.02 1.205 5.02 1.145 4.67 1.145 4.67 1.205 4.61 1.205 4.61 1.145 4.26 1.145 4.26 1.205 4.2 1.205 4.2 1.145 3.85 1.145 3.85 1.205 3.79 1.205 3.79 1.145 3.44 1.145 3.44 1.205 3.38 1.205 3.38 1.055 3.03 1.055 3.03 1.115 2.97 1.115 2.97 0.895 2.74 0.895 2.74 0.92 2.64 0.92 2.64 0.395 0.955 0.395 0.955 0.335 4.6 0.335 4.6 0.395 2.7 0.395 2.7 0.79 2.74 0.79 2.74 0.815 3.03 0.815 3.03 0.995 3.44 0.995 3.44 1.085 5.08 1.085 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.69230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.165 0.895 2.125 0.895 2.125 0.935 2.095 0.935 2.095 0.985 1.23 0.985 1.23 0.905 0.975 0.905 0.975 0.845 1.29 0.845 1.29 0.925 2.035 0.925 2.035 0.815 2.165 0.815 ;
    END
  END A2
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.576923 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.57 0.895 4.34 0.895 4.34 0.985 3.54 0.985 3.54 0.895 3.435 0.895 3.435 0.815 3.6 0.815 3.6 0.925 4.28 0.925 4.28 0.835 4.57 0.835 ;
    END
  END B2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.9615385 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.95 0.895 4.94 0.895 4.94 0.92 4.86 0.92 4.86 0.835 4.67 0.835 4.67 0.735 4.18 0.735 4.18 0.825 3.7 0.825 3.7 0.715 3.07 0.715 3.07 0.655 3.76 0.655 3.76 0.765 4.12 0.765 4.12 0.675 4.73 0.675 4.73 0.775 4.95 0.775 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.602564 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.36 0.715 1.935 0.715 1.935 0.825 1.39 0.825 1.39 0.745 0.74 0.745 0.74 0.92 0.66 0.92 0.66 0.85 0.6 0.85 0.6 0.79 0.68 0.79 0.68 0.685 1.45 0.685 1.45 0.765 1.875 0.765 1.875 0.655 2.36 0.655 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.62820525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.54 0.73 2.46 0.73 2.46 0.555 1.67 0.555 1.67 0.665 1.55 0.665 1.55 0.555 0.5 0.555 0.5 0.695 0.44 0.695 0.44 0.495 2.54 0.495 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.025641 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.11 0.705 5.05 0.705 5.05 0.555 4.02 0.555 4.02 0.665 3.9 0.665 3.9 0.555 2.965 0.555 2.965 0.665 2.8 0.665 2.8 0.585 2.905 0.585 2.905 0.495 5.11 0.495 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 1.77 0 1.77 0 1.65 0.455 1.65 0.455 1.245 0.515 1.245 0.515 1.65 0.865 1.65 0.865 1.245 0.925 1.245 0.925 1.65 1.295 1.65 1.295 1.245 1.355 1.245 1.355 1.65 1.72 1.65 1.72 1.245 1.78 1.245 1.78 1.65 2.13 1.65 2.13 1.245 2.19 1.245 2.19 1.65 2.54 1.65 2.54 1.245 2.6 1.245 2.6 1.65 5.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 0.06 5.155 0.06 5.155 0.305 5.215 0.305 5.215 0.365 5.095 0.365 5.095 0.06 4.1 0.06 4.1 0.17 3.98 0.17 3.98 0.06 2.765 0.06 2.765 0.17 2.645 0.17 2.645 0.06 1.575 0.06 1.575 0.17 1.455 0.17 1.455 0.06 0.425 0.06 0.425 0.305 0.485 0.305 0.485 0.365 0.365 0.365 0.365 0.06 0 0.06 0 -0.06 5.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.285 1.365 2.745 1.365 2.745 1.145 2.395 1.145 2.395 1.365 2.335 1.365 2.335 1.145 1.985 1.145 1.985 1.365 1.925 1.365 1.925 1.145 1.575 1.145 1.575 1.365 1.515 1.365 1.515 1.145 1.13 1.145 1.13 1.365 1.07 1.365 1.07 1.145 0.72 1.145 0.72 1.365 0.66 1.365 0.66 1.08 0.31 1.08 0.31 1.365 0.25 1.365 0.25 0.975 0.31 0.975 0.31 1.02 0.72 1.02 0.72 1.085 1.07 1.085 1.07 1.005 1.13 1.005 1.13 1.085 2.335 1.085 2.335 0.975 2.395 0.975 2.395 1.085 2.745 1.085 2.745 1.02 2.805 1.02 2.805 1.305 3.175 1.305 3.175 1.245 3.235 1.245 3.235 1.305 3.585 1.305 3.585 1.245 3.645 1.245 3.645 1.305 3.995 1.305 3.995 1.245 4.055 1.245 4.055 1.305 4.405 1.305 4.405 1.245 4.465 1.245 4.465 1.305 4.815 1.305 4.815 1.245 4.875 1.245 4.875 1.305 5.225 1.305 5.225 0.975 5.285 0.975 ;
  END
END AOI33X4

MACRO AOI33XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI33XL 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5895 LAYER Metal1 ;
    ANTENNADIFFAREA 0.7605 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.35 1.3 1.26 1.3 1.26 1.17 0.91 1.17 0.91 1.265 0.85 1.265 0.85 1.11 1.26 1.11 1.26 0.41 0.645 0.41 0.645 0.29 0.705 0.29 0.705 0.35 1.32 0.35 1.32 1.17 1.35 1.17 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.12962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.26 1.11 0.06 1.11 0.06 0.925 0.165 0.925 0.165 0.995 0.26 0.995 ;
    END
  END A0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.388889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.595 0.66 0.74 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.64814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.97 0.63 0.95 0.63 0.95 0.975 0.86 0.975 0.86 0.51 0.97 0.51 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.51 1.15 1.01 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.47 0.895 0.4 0.895 0.4 0.92 0.26 0.92 0.26 0.765 0.375 0.765 0.375 0.805 0.47 0.805 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.92 0.78 1.11 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.08 1.65 0.08 1.51 0.14 1.51 0.14 1.65 0.41 1.65 0.41 1.51 0.47 1.51 0.47 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 1.225 0.06 1.225 0.19 1.285 0.19 1.285 0.25 1.165 0.25 1.165 0.06 0.165 0.06 0.165 0.41 0.105 0.41 0.105 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.145 1.33 1.07 1.33 1.07 1.425 0.645 1.425 0.645 1.3 0.215 1.3 0.215 1.24 0.705 1.24 0.705 1.365 1.01 1.365 1.01 1.27 1.145 1.27 ;
  END
END AOI33XL

MACRO BMXIX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BMXIX2 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN PPN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3124 LAYER Metal1 ;
    ANTENNADIFFAREA 2.487425 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1071 LAYER Metal1 ;
      ANTENNAMAXAREACAR 21.5910365 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 169.439776 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.06 0.54 4.14 1.29 ;
    END
  END PPN
  PIN X2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.525 3.74 1.025 ;
    END
  END X2
  PIN M1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.78 0.815 2.28 0.895 ;
    END
  END M1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.44 0.895 1.315 0.895 1.315 0.96 1.165 0.96 1.165 0.88 1.235 0.88 1.235 0.655 1.44 0.655 ;
    END
  END A
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 18.6574075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.005 1.44 0.57 1.44 0.57 1.095 0.505 1.095 0.505 1.085 0.435 1.085 0.435 1.005 0.445 1.005 0.445 0.995 0.565 0.995 0.565 1.035 0.63 1.035 0.63 1.38 2.005 1.38 ;
    END
  END S
  PIN M0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.745 0.935 0.665 0.935 0.665 0.895 0.33 0.895 0.33 0.935 0.25 0.935 0.25 0.895 0.235 0.895 0.235 0.815 0.745 0.815 ;
    END
  END M0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.41 1.65 0.41 1.22 0.47 1.22 0.47 1.65 1.185 1.65 1.185 1.54 1.305 1.54 1.305 1.65 2.065 1.65 2.065 1.54 2.185 1.54 2.185 1.65 3.82 1.65 3.82 1.095 3.88 1.095 3.88 1.65 4.265 1.65 4.265 0.9 4.325 0.9 4.325 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 4.325 0.06 4.325 0.52 4.265 0.52 4.265 0.06 3.915 0.06 3.915 0.17 3.795 0.17 3.795 0.06 2.185 0.06 2.185 0.17 2.065 0.17 2.065 0.06 1.225 0.06 1.225 0.555 1.165 0.555 1.165 0.06 0.395 0.06 0.395 0.555 0.335 0.555 0.335 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.96 0.82 3.9 0.82 3.9 0.425 3.635 0.425 3.635 0.415 3.125 0.415 3.125 1.145 3.065 1.145 3.065 0.355 3.695 0.355 3.695 0.365 3.96 0.365 ;
      POLYGON 3.705 1.185 3.49 1.185 3.49 1.465 2.995 1.465 2.995 1.405 3.43 1.405 3.43 0.735 3.44 0.735 3.44 0.57 3.56 0.57 3.56 0.63 3.5 0.63 3.5 0.795 3.49 0.795 3.49 1.125 3.705 1.125 ;
      POLYGON 3.33 1.305 2.895 1.305 2.895 1.375 2.105 1.375 2.105 1.28 1.64 1.28 1.64 1.22 2.165 1.22 2.165 1.315 2.835 1.315 2.835 1.245 2.905 1.245 2.905 0.395 1.815 0.395 1.815 0.555 1.755 0.555 1.755 0.335 2.965 0.335 2.965 1.245 3.27 1.245 3.27 0.515 3.33 0.515 ;
      POLYGON 2.805 0.66 2.735 0.66 2.735 1.025 2.805 1.025 2.805 1.145 2.735 1.145 2.735 1.215 2.265 1.215 2.265 1.12 0.905 1.12 0.905 1.215 0.785 1.215 0.785 1.155 0.845 1.155 0.845 0.55 0.655 0.55 0.655 0.49 0.905 0.49 0.905 1.06 2.325 1.06 2.325 1.155 2.675 1.155 2.675 0.6 2.745 0.6 2.745 0.54 2.805 0.54 ;
      POLYGON 2.545 1.055 2.425 1.055 2.425 0.995 2.485 0.995 2.485 0.715 1.6 0.715 1.6 0.885 1.54 0.885 1.54 0.655 2.485 0.655 2.485 0.555 2.3 0.555 2.3 0.495 2.545 0.495 ;
      POLYGON 1.065 0.885 1.005 0.885 1.005 0.39 0.555 0.39 0.555 0.655 0.67 0.655 0.67 0.715 0.135 0.715 0.135 1.035 0.265 1.035 0.265 1.245 0.205 1.245 0.205 1.095 0.075 1.095 0.075 0.655 0.13 0.655 0.13 0.46 0.19 0.46 0.19 0.655 0.495 0.655 0.495 0.33 1.065 0.33 ;
  END
END BMXIX2

MACRO BMXIX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BMXIX4 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN M1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 15.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.405 0.855 1.815 0.855 1.815 0.25 1.59 0.25 1.59 0.19 1.53 0.19 1.53 0.13 1.65 0.13 1.65 0.19 1.875 0.19 1.875 0.625 1.965 0.625 1.965 0.795 2.345 0.795 2.345 0.735 2.405 0.735 ;
    END
  END M1
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.45 1.34 0.95 ;
    END
  END A
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 20.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.085 1.335 1.06 1.335 1.06 1.27 0.66 1.27 0.66 0.82 0.4 0.82 0.4 0.76 0.72 0.76 0.72 0.98 0.74 0.98 0.74 1.21 1.12 1.21 1.12 1.275 2.085 1.275 ;
    END
  END S
  PIN M0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 12.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.96 1.43 0.5 1.43 0.5 1.275 0.235 1.275 0.235 0.765 0.295 0.765 0.295 1.195 0.365 1.195 0.365 1.215 0.56 1.215 0.56 1.37 0.96 1.37 ;
    END
  END M0
  PIN PPN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.52805 LAYER Metal1 ;
    ANTENNADIFFAREA 3.0339 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.17865 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.1508535 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 107.22082275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.725 1.29 4.665 1.29 4.665 0.73 4.315 0.73 4.315 1.29 4.255 1.29 4.255 0.54 4.315 0.54 4.315 0.6 4.34 0.6 4.34 0.67 4.665 0.67 4.665 0.54 4.725 0.54 ;
    END
  END PPN
  PIN X2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.05280525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.565 1.465 3.435 1.465 3.435 1.445 3.165 1.445 3.165 0.855 3.075 0.855 3.075 0.735 3.225 0.735 3.225 1.385 3.565 1.385 ;
    END
  END X2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 1.77 0 1.77 0 1.65 0.3 1.65 0.3 1.54 0.42 1.54 0.42 1.65 1.255 1.65 1.255 1.54 1.375 1.54 1.375 1.65 2.135 1.65 2.135 1.54 2.255 1.54 2.255 1.65 4.02 1.65 4.02 1.285 4.08 1.285 4.08 1.65 4.46 1.65 4.46 0.9 4.52 0.9 4.52 1.65 4.87 1.65 4.87 0.9 4.93 0.9 4.93 1.65 5 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 0.06 4.93 0.06 4.93 0.52 4.87 0.52 4.87 0.06 4.52 0.06 4.52 0.52 4.46 0.52 4.46 0.06 4.11 0.06 4.11 0.635 4.05 0.635 4.05 0.06 2.4 0.06 2.4 0.2 2.34 0.2 2.34 0.06 1.29 0.06 1.29 0.35 1.17 0.35 1.17 0.06 0.36 0.06 0.36 0.38 0.3 0.38 0.3 0.06 0 0.06 0 -0.06 5 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.155 1.185 3.92 1.185 3.92 1.2 3.325 1.2 3.325 0.63 3.09 0.63 3.09 0.55 3.21 0.55 3.21 0.57 3.385 0.57 3.385 1.14 3.86 1.14 3.86 1.125 4.095 1.125 4.095 0.74 4.155 0.74 ;
      POLYGON 3.905 1.02 3.825 1.02 3.825 0.74 3.645 0.74 3.645 0.66 3.825 0.66 3.825 0.54 3.905 0.54 ;
      POLYGON 3.59 1.04 3.53 1.04 3.53 0.98 3.485 0.98 3.485 0.47 3.31 0.47 3.31 0.42 2.815 0.42 2.815 1.175 2.345 1.175 2.345 1.015 1.655 1.015 1.655 0.375 1.595 0.375 1.595 0.315 1.715 0.315 1.715 0.955 2.405 0.955 2.405 1.115 2.755 1.115 2.755 0.36 3.37 0.36 3.37 0.41 3.545 0.41 3.545 0.92 3.59 0.92 ;
      POLYGON 3.065 1.335 2.185 1.335 2.185 1.175 1.22 1.175 1.22 1.11 0.85 1.11 0.85 0.375 0.71 0.375 0.71 0.315 0.91 0.315 0.91 1.05 1.28 1.05 1.28 1.115 2.245 1.115 2.245 1.275 3.005 1.275 3.005 1.015 2.915 1.015 2.915 0.52 2.975 0.52 2.975 0.955 3.065 0.955 ;
      POLYGON 2.625 1.015 2.505 1.015 2.505 0.635 2.125 0.635 2.125 0.695 2.065 0.695 2.065 0.575 2.505 0.575 2.505 0.515 2.565 0.515 2.565 0.955 2.625 0.955 ;
      POLYGON 1.07 0.885 1.01 0.885 1.01 0.22 0.61 0.22 0.61 0.51 0.75 0.51 0.75 0.57 0.135 0.57 0.135 1.045 0.075 1.045 0.075 0.285 0.135 0.285 0.135 0.51 0.55 0.51 0.55 0.16 1.07 0.16 ;
  END
END BMXIX4

MACRO BUFX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX12 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.89745 LAYER Metal1 ;
    ANTENNADIFFAREA 2.3684 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.351 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.4058405 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 43.905983 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.98 0.655 0.295 0.655 0.295 0.98 1.98 0.98 1.98 1.45 1.92 1.45 1.92 1.04 1.57 1.04 1.57 1.45 1.51 1.45 1.51 1.04 1.16 1.04 1.16 1.45 1.1 1.45 1.1 1.04 0.75 1.04 0.75 1.45 0.69 1.45 0.69 1.04 0.34 1.04 0.34 1.45 0.26 1.45 0.26 1.04 0.215 1.04 0.215 0.595 0.28 0.595 0.28 0.255 0.34 0.255 0.34 0.595 0.69 0.595 0.69 0.255 0.75 0.255 0.75 0.595 1.1 0.595 1.1 0.255 1.16 0.255 1.16 0.595 1.51 0.595 1.51 0.255 1.57 0.255 1.57 0.595 1.92 0.595 1.92 0.255 1.98 0.255 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.08775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.17948725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.45 0.795 2.715 0.875 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.77 0 1.77 0 1.65 0.075 1.65 0.075 0.98 0.135 0.98 0.135 1.65 0.485 1.65 0.485 1.14 0.545 1.14 0.545 1.65 0.895 1.65 0.895 1.14 0.955 1.14 0.955 1.65 1.305 1.65 1.305 1.14 1.365 1.14 1.365 1.65 1.715 1.65 1.715 1.14 1.775 1.14 1.775 1.65 2.125 1.65 2.125 1.14 2.185 1.14 2.185 1.65 2.535 1.65 2.535 1.14 2.595 1.14 2.595 1.65 3 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 0.06 2.595 0.06 2.595 0.565 2.535 0.565 2.535 0.06 2.185 0.06 2.185 0.565 2.125 0.565 2.125 0.06 1.775 0.06 1.775 0.53 1.715 0.53 1.715 0.06 1.365 0.06 1.365 0.53 1.305 0.53 1.305 0.06 0.955 0.06 0.955 0.53 0.895 0.53 0.895 0.06 0.545 0.06 0.545 0.53 0.485 0.53 0.485 0.06 0.135 0.06 0.135 0.565 0.075 0.565 0.075 0.06 0 0.06 0 -0.06 3 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.8 0.695 2.39 0.695 2.39 1 2.8 1 2.8 1.45 2.74 1.45 2.74 1.065 2.39 1.065 2.39 1.45 2.33 1.45 2.33 0.785 0.395 0.785 0.395 0.725 2.33 0.725 2.33 0.305 2.39 0.305 2.39 0.635 2.74 0.635 2.74 0.305 2.8 0.305 ;
  END
END BUFX12

MACRO BUFX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX16 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.553675 LAYER Metal1 ;
    ANTENNADIFFAREA 3.2877 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4662 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.47763825 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 44.20205925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.795 0.685 0.315 0.685 0.315 0.905 2.795 0.905 2.795 1.345 2.735 1.345 2.735 0.965 2.385 0.965 2.385 1.345 2.325 1.345 2.325 0.965 1.975 0.965 1.975 1.345 1.915 1.345 1.915 0.965 1.565 0.965 1.565 1.345 1.505 1.345 1.505 0.965 1.155 0.965 1.155 1.345 1.095 1.345 1.095 0.965 0.745 0.965 0.745 1.345 0.685 1.345 0.685 0.965 0.335 0.965 0.335 1.345 0.235 1.345 0.235 0.365 0.335 0.365 0.335 0.625 0.685 0.625 0.685 0.365 0.745 0.365 0.745 0.625 1.095 0.625 1.095 0.365 1.155 0.365 1.155 0.625 1.505 0.625 1.505 0.365 1.565 0.365 1.565 0.625 1.915 0.625 1.915 0.365 1.975 0.365 1.975 0.625 2.325 0.625 2.325 0.365 2.385 0.365 2.385 0.625 2.735 0.625 2.735 0.365 2.795 0.365 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.64102575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.265 0.755 3.825 0.835 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.9 0.13 0.9 0.13 1.65 0.48 1.65 0.48 1.065 0.54 1.065 0.54 1.65 0.89 1.65 0.89 1.065 0.95 1.065 0.95 1.65 1.3 1.65 1.3 1.065 1.36 1.065 1.36 1.65 1.71 1.65 1.71 1.065 1.77 1.065 1.77 1.65 2.12 1.65 2.12 1.065 2.18 1.065 2.18 1.65 2.53 1.65 2.53 1.065 2.59 1.065 2.59 1.65 2.94 1.65 2.94 0.955 3 0.955 3 1.65 3.35 1.65 3.35 1.07 3.41 1.07 3.41 1.65 3.76 1.65 3.76 0.955 3.82 0.955 3.82 1.65 4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.82 0.06 3.82 0.66 3.76 0.66 3.76 0.06 3.41 0.06 3.41 0.52 3.35 0.52 3.35 0.06 3 0.06 3 0.66 2.94 0.66 2.94 0.06 2.59 0.06 2.59 0.485 2.53 0.485 2.53 0.06 2.18 0.06 2.18 0.485 2.12 0.485 2.12 0.06 1.77 0.06 1.77 0.485 1.71 0.485 1.71 0.06 1.36 0.06 1.36 0.485 1.3 0.485 1.3 0.06 0.95 0.06 0.95 0.485 0.89 0.485 0.89 0.06 0.54 0.06 0.54 0.485 0.48 0.485 0.48 0.06 0.13 0.06 0.13 0.66 0.07 0.66 0.07 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.615 0.68 3.205 0.68 3.205 0.73 3.185 0.73 3.185 0.86 3.205 0.86 3.205 0.895 3.615 0.895 3.615 1.345 3.555 1.345 3.555 0.955 3.205 0.955 3.205 1.345 3.145 1.345 3.145 0.925 3.11 0.925 3.11 0.805 0.395 0.805 0.395 0.745 3.11 0.745 3.11 0.66 3.145 0.66 3.145 0.4 3.205 0.4 3.205 0.62 3.555 0.62 3.555 0.4 3.615 0.4 ;
  END
END BUFX16

MACRO BUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX2 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4539 LAYER Metal1 ;
    ANTENNADIFFAREA 0.572 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.75897425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 65.74358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.335 1.32 0.275 1.32 0.275 0.88 0.185 0.88 0.185 0.76 0.275 0.76 0.275 0.38 0.335 0.38 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.5555555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.565 0.76 0.745 0.88 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.93 0.13 0.93 0.13 1.65 0.48 1.65 0.48 1.185 0.54 1.185 0.54 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.54 0.06 0.54 0.5 0.48 0.5 0.48 0.06 0.13 0.06 0.13 0.64 0.07 0.64 0.07 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.745 0.7 0.48 0.7 0.48 0.94 0.745 0.94 0.745 1.235 0.685 1.235 0.685 1 0.42 1 0.42 0.64 0.685 0.64 0.685 0.405 0.745 0.405 ;
  END
END BUFX2

MACRO BUFX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX20 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.10005 LAYER Metal1 ;
    ANTENNADIFFAREA 3.84 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.585225 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.2971935 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 43.291042 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.41 0.715 0.14 0.715 0.14 0.92 3.41 0.92 3.41 1.365 3.35 1.365 3.35 0.98 3 0.98 3 1.365 2.94 1.365 2.94 0.98 2.59 0.98 2.59 1.365 2.53 1.365 2.53 0.98 2.18 0.98 2.18 1.365 2.12 1.365 2.12 0.98 1.77 0.98 1.77 1.365 1.71 1.365 1.71 0.98 1.36 0.98 1.36 1.365 1.3 1.365 1.3 0.98 0.95 0.98 0.95 1.365 0.89 1.365 0.89 0.98 0.54 0.98 0.54 1.365 0.48 1.365 0.48 0.98 0.13 0.98 0.13 1.365 0.06 1.365 0.06 0.355 0.13 0.355 0.13 0.655 0.48 0.655 0.48 0.355 0.54 0.355 0.54 0.655 0.89 0.655 0.89 0.355 0.95 0.355 0.95 0.655 1.3 0.655 1.3 0.355 1.36 0.355 1.36 0.655 1.71 0.655 1.71 0.355 1.77 0.355 1.77 0.655 2.12 0.655 2.12 0.355 2.18 0.355 2.18 0.655 2.53 0.655 2.53 0.355 2.59 0.355 2.59 0.655 2.94 0.655 2.94 0.355 3 0.355 3 0.655 3.35 0.655 3.35 0.355 3.41 0.355 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.14625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.1897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.875 0.76 4.375 0.84 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.08 0.335 1.08 0.335 1.65 0.685 1.65 0.685 1.08 0.745 1.08 0.745 1.65 1.095 1.65 1.095 1.08 1.155 1.08 1.155 1.65 1.505 1.65 1.505 1.08 1.565 1.08 1.565 1.65 1.915 1.65 1.915 1.08 1.975 1.08 1.975 1.65 2.325 1.65 2.325 1.08 2.385 1.08 2.385 1.65 2.735 1.65 2.735 1.08 2.795 1.08 2.795 1.65 3.145 1.65 3.145 1.08 3.205 1.08 3.205 1.65 3.555 1.65 3.555 0.975 3.615 0.975 3.615 1.65 3.965 1.65 3.965 1.125 4.025 1.125 4.025 1.65 4.375 1.65 4.375 1.125 4.435 1.125 4.435 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 4.435 0.06 4.435 0.52 4.375 0.52 4.375 0.06 4.025 0.06 4.025 0.52 3.965 0.52 3.965 0.06 3.615 0.06 3.615 0.64 3.555 0.64 3.555 0.06 3.205 0.06 3.205 0.595 3.145 0.595 3.145 0.06 2.795 0.06 2.795 0.595 2.735 0.595 2.735 0.06 2.385 0.06 2.385 0.595 2.325 0.595 2.325 0.06 1.975 0.06 1.975 0.595 1.915 0.595 1.915 0.06 1.565 0.06 1.565 0.595 1.505 0.595 1.505 0.06 1.155 0.06 1.155 0.595 1.095 0.595 1.095 0.06 0.745 0.06 0.745 0.595 0.685 0.595 0.685 0.06 0.335 0.06 0.335 0.595 0.275 0.595 0.275 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.64 0.68 3.775 0.68 3.775 1 4.64 1 4.64 1.365 4.58 1.365 4.58 1.06 4.23 1.06 4.23 1.365 4.17 1.365 4.17 1.06 3.82 1.06 3.82 1.365 3.76 1.365 3.76 1.06 3.715 1.06 3.715 0.835 0.31 0.835 0.31 0.775 3.715 0.775 3.715 0.62 3.76 0.62 3.76 0.4 3.82 0.4 3.82 0.62 4.17 0.62 4.17 0.4 4.23 0.4 4.23 0.62 4.58 0.62 4.58 0.4 4.64 0.4 ;
  END
END BUFX20

MACRO BUFX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX3 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6685 LAYER Metal1 ;
    ANTENNADIFFAREA 0.782 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.08775 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.6182335 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 62.18803425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 1.44 0.48 1.44 0.48 0.955 0.13 0.955 0.13 1.44 0.07 1.44 0.07 0.86 0.05 0.86 0.05 0.78 0.07 0.78 0.07 0.34 0.13 0.34 0.13 0.895 0.48 0.895 0.48 0.345 0.54 0.345 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.945 0.86 0.76 0.86 0.76 0.73 0.925 0.73 0.925 0.78 0.945 0.78 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.05 0.335 1.05 0.335 1.65 0.685 1.65 0.685 1.08 0.745 1.08 0.745 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.745 0.06 0.745 0.51 0.685 0.51 0.685 0.06 0.335 0.06 0.335 0.6 0.275 0.6 0.275 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.95 0.67 0.695 0.67 0.695 0.96 0.95 0.96 0.95 1.44 0.89 1.44 0.89 1.02 0.635 1.02 0.635 0.61 0.89 0.61 0.89 0.34 0.95 0.34 ;
  END
END BUFX3

MACRO BUFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX4 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8055 LAYER Metal1 ;
    ANTENNADIFFAREA 0.94375 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.8846155 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 55.25641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 1.37 0.7 1.37 0.7 0.86 0.335 0.86 0.335 1.37 0.275 1.37 0.275 0.86 0.07 0.86 0.07 0.78 0.275 0.78 0.275 0.23 0.335 0.23 0.335 0.78 0.7 0.78 0.7 0.23 0.76 0.23 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5384615 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.17 0.86 1.145 0.86 1.145 0.91 1.015 0.91 1.015 0.72 1.145 0.72 1.145 0.78 1.17 0.78 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.98 0.13 0.98 0.13 1.65 0.48 1.65 0.48 0.98 0.54 0.98 0.54 1.65 0.905 1.65 0.905 1.115 0.965 1.115 0.965 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 0.965 0.06 0.965 0.48 0.905 0.48 0.905 0.06 0.54 0.06 0.54 0.48 0.48 0.48 0.48 0.06 0.13 0.06 0.13 0.48 0.07 0.48 0.07 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.17 0.66 0.945 0.66 0.945 0.97 1.17 0.97 1.17 1.37 1.11 1.37 1.11 1.03 0.885 1.03 0.885 0.66 0.825 0.66 0.825 0.6 1.11 0.6 1.11 0.23 1.17 0.23 ;
  END
END BUFX4

MACRO BUFX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX6 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.565 0.06 1.565 0.59 1.505 0.59 1.505 0.06 1.155 0.06 1.155 0.61 1.095 0.61 1.095 0.06 0.745 0.06 0.745 0.625 0.685 0.625 0.685 0.06 0.335 0.06 0.335 0.625 0.275 0.625 0.275 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.275 1.65 0.275 0.985 0.335 0.985 0.335 1.65 0.685 1.65 0.685 0.985 0.745 0.985 0.745 1.65 1.095 1.65 1.095 0.915 1.155 0.915 1.155 1.65 1.505 1.65 1.505 0.9 1.565 0.9 1.565 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.6153845 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.425 0.665 1.565 0.84 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.04355 LAYER Metal1 ;
    ANTENNADIFFAREA 1.3524 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.94615375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 47.79487175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.95 1.37 0.89 1.37 0.89 0.895 0.54 0.895 0.54 1.37 0.48 1.37 0.48 0.895 0.13 0.895 0.13 1.37 0.06 1.37 0.06 0.35 0.13 0.35 0.13 0.76 0.14 0.76 0.14 0.835 0.48 0.835 0.48 0.35 0.54 0.35 0.54 0.835 0.89 0.835 0.89 0.35 0.95 0.35 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      POLYGON 1.36 1.29 1.3 1.29 1.3 0.805 1.015 0.805 1.015 0.745 1.3 0.745 1.3 0.35 1.36 0.35 ;
  END
END BUFX6

MACRO BUFX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX8 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3243 LAYER Metal1 ;
    ANTENNADIFFAREA 1.65 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.68125275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 46.3963965 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.515 0.705 0.285 0.705 0.285 0.93 1.515 0.93 1.515 1.375 1.455 1.375 1.455 0.99 1.105 0.99 1.105 1.375 1.045 1.375 1.045 0.99 0.695 0.99 0.695 1.375 0.635 1.375 0.635 0.99 0.285 0.99 0.285 1.375 0.225 1.375 0.225 0.84 0.205 0.84 0.205 0.76 0.225 0.76 0.225 0.345 0.285 0.345 0.285 0.645 0.635 0.645 0.635 0.345 0.695 0.345 0.695 0.645 1.045 0.645 1.045 0.345 1.105 0.345 1.105 0.645 1.455 0.645 1.455 0.345 1.515 0.345 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.69230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.16 0.845 2 0.845 2 0.675 2.15 0.675 2.15 0.765 2.16 0.765 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.43 1.65 0.43 1.09 0.49 1.09 0.49 1.65 0.84 1.65 0.84 1.09 0.9 1.09 0.9 1.65 1.25 1.65 1.25 1.09 1.31 1.09 1.31 1.65 1.66 1.65 1.66 0.93 1.72 0.93 1.72 1.65 2.07 1.65 2.07 0.93 2.13 0.93 2.13 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 2.13 0.06 2.13 0.5 2.07 0.5 2.07 0.06 1.72 0.06 1.72 0.5 1.66 0.5 1.66 0.06 1.31 0.06 1.31 0.585 1.25 0.585 1.25 0.06 0.9 0.06 0.9 0.585 0.84 0.585 0.84 0.06 0.49 0.06 0.49 0.585 0.43 0.585 0.43 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.925 1.32 1.865 1.32 1.865 0.825 0.54 0.825 0.54 0.765 1.865 0.765 1.865 0.52 1.925 0.52 ;
  END
END BUFX8

MACRO CLKAND2X12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X12 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.357575 LAYER Metal1 ;
    ANTENNADIFFAREA 3.38565 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.351 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.716738 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 52.16239325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.14 1.37 4.035 1.37 4.035 0.975 3.685 0.975 3.685 1.37 3.625 1.37 3.625 0.975 3.275 0.975 3.275 1.37 3.215 1.37 3.215 0.975 2.865 0.975 2.865 1.37 2.805 1.37 2.805 0.975 2.455 0.975 2.455 1.37 2.395 1.37 2.395 0.915 4.06 0.915 4.06 0.655 2.305 0.655 2.305 0.35 2.365 0.35 2.365 0.595 2.715 0.595 2.715 0.35 2.775 0.35 2.775 0.595 3.125 0.595 3.125 0.35 3.185 0.35 3.185 0.595 3.535 0.595 3.535 0.35 3.595 0.35 3.595 0.595 3.945 0.595 3.945 0.35 4.005 0.35 4.005 0.595 4.12 0.595 4.12 0.79 4.14 0.79 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.122625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.1590215 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.045 0.875 1.965 0.875 1.965 1.01 0.66 1.01 0.66 0.89 0.72 0.89 0.72 0.95 1.19 0.95 1.19 0.89 1.25 0.89 1.25 0.95 1.835 0.95 1.835 0.815 2.045 0.815 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.122625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.64 0.85 1.58 0.85 1.58 0.79 1.085 0.79 1.085 0.8 0.965 0.8 0.965 0.79 0.54 0.79 0.54 0.92 0.46 0.92 0.46 0.85 0.265 0.85 0.265 0.79 0.48 0.79 0.48 0.73 1.64 0.73 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.12 1.65 0.12 1.165 0.18 1.165 0.18 1.65 0.56 1.65 0.56 1.51 0.62 1.51 0.62 1.65 0.96 1.65 0.96 1.51 1.02 1.51 1.02 1.65 1.36 1.65 1.36 1.51 1.42 1.51 1.42 1.65 1.76 1.65 1.76 1.51 1.82 1.51 1.82 1.65 2.16 1.65 2.16 1.51 2.22 1.51 2.22 1.65 2.6 1.65 2.6 1.075 2.66 1.075 2.66 1.65 3.01 1.65 3.01 1.075 3.07 1.075 3.07 1.65 3.42 1.65 3.42 1.075 3.48 1.075 3.48 1.65 3.83 1.65 3.83 1.075 3.89 1.075 3.89 1.65 4.24 1.65 4.24 0.9 4.3 0.9 4.3 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 4.28 0.06 4.28 0.66 4.22 0.66 4.22 0.06 3.8 0.06 3.8 0.47 3.74 0.47 3.74 0.06 3.39 0.06 3.39 0.47 3.33 0.47 3.33 0.06 2.98 0.06 2.98 0.47 2.92 0.47 2.92 0.06 2.57 0.06 2.57 0.47 2.51 0.47 2.51 0.06 2.09 0.06 2.09 0.47 2.03 0.47 2.03 0.06 1.315 0.06 1.315 0.47 1.255 0.47 1.255 0.06 0.615 0.06 0.615 0.47 0.555 0.47 0.555 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.96 0.815 2.205 0.815 2.205 1.17 0.295 1.17 0.295 1.11 2.145 1.11 2.145 0.63 0.22 0.63 0.22 0.35 0.28 0.35 0.28 0.57 0.865 0.57 0.865 0.51 0.925 0.51 0.925 0.57 1.72 0.57 1.72 0.35 1.78 0.35 1.78 0.57 2.205 0.57 2.205 0.755 3.96 0.755 ;
  END
END CLKAND2X12

MACRO CLKAND2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X2 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5735 LAYER Metal1 ;
    ANTENNADIFFAREA 0.763225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.80341875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 76.15384625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 0.73 0.86 0.73 0.86 0.88 0.765 0.88 0.765 1.34 0.705 1.34 0.705 0.82 0.8 0.82 0.8 0.42 0.705 0.42 0.705 0.3 0.765 0.3 0.765 0.36 0.86 0.36 0.86 0.6 0.94 0.6 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.022725 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.65676575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 1.12 0.46 1.12 0.46 1.06 0.4 1.06 0.4 0.68 0.485 0.68 0.485 0.98 0.54 0.98 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.022725 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.65676575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.79 0.14 1.29 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.08 1.65 0.08 1.51 0.14 1.51 0.14 1.65 0.5 1.65 0.5 1.22 0.56 1.22 0.56 1.65 0.96 1.65 0.96 0.95 1.02 0.95 1.02 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 1.02 0.06 1.02 0.42 0.96 0.42 0.96 0.06 0.56 0.06 0.56 0.42 0.5 0.42 0.5 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.7 0.72 0.64 0.72 0.64 0.58 0.3 0.58 0.3 1.245 0.24 1.245 0.24 0.56 0.16 0.56 0.16 0.5 0.3 0.5 0.3 0.52 0.7 0.52 ;
  END
END CLKAND2X2

MACRO CLKAND2X3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X3 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8362 LAYER Metal1 ;
    ANTENNADIFFAREA 1.15195 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.08775 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.52934475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 72.13675225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.625 1.335 1.565 1.335 1.565 1.005 1.215 1.005 1.215 1.335 1.155 1.335 1.155 0.945 1.46 0.945 1.46 0.555 1.125 0.555 1.125 0.505 1.065 0.505 1.065 0.445 1.185 0.445 1.185 0.495 1.505 0.495 1.505 0.415 1.565 0.415 1.565 0.555 1.54 0.555 1.54 0.945 1.625 0.945 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04095 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.36996325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.805 0.57 0.925 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04095 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.908425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.215 0.625 0.805 0.705 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.02 0.13 1.02 0.13 1.65 0.51 1.65 0.51 1.51 0.57 1.51 0.57 1.65 0.92 1.65 0.92 1.51 0.98 1.51 0.98 1.65 1.36 1.65 1.36 1.105 1.42 1.105 1.42 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.36 0.06 1.36 0.395 1.3 0.395 1.3 0.06 0.82 0.06 0.82 0.305 0.88 0.305 0.88 0.365 0.76 0.365 0.76 0.06 0.23 0.06 0.23 0.395 0.17 0.395 0.17 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.18 0.715 0.965 0.715 0.965 1.085 0.245 1.085 0.245 1.025 0.905 1.025 0.905 0.525 0.52 0.525 0.52 0.505 0.45 0.505 0.45 0.445 0.57 0.445 0.57 0.465 0.965 0.465 0.965 0.655 1.18 0.655 ;
  END
END CLKAND2X3

MACRO CLKAND2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X4 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.95105 LAYER Metal1 ;
    ANTENNADIFFAREA 1.3256 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.1286325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 61.3846155 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 1.335 1.645 1.335 1.645 1.005 1.295 1.005 1.295 1.335 1.235 1.335 1.235 0.945 1.66 0.945 1.66 0.565 1.135 0.565 1.135 0.425 1.195 0.425 1.195 0.505 1.545 0.505 1.545 0.425 1.605 0.425 1.605 0.505 1.72 0.505 1.72 0.79 1.74 0.79 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04095 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.24908425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.265 0.815 0.765 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04095 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.981685 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.875 0.715 0.285 0.715 0.285 0.635 0.435 0.635 0.435 0.625 0.565 0.625 0.565 0.635 0.875 0.635 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.18 1.65 0.18 1.51 0.24 1.51 0.24 1.65 0.51 1.65 0.51 1.51 0.57 1.51 0.57 1.65 1 1.65 1 1.51 1.06 1.51 1.06 1.65 1.44 1.65 1.44 1.105 1.5 1.105 1.5 1.65 1.85 1.65 1.85 0.945 1.91 0.945 1.91 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.81 0.06 1.81 0.405 1.75 0.405 1.75 0.06 1.4 0.06 1.4 0.405 1.34 0.405 1.34 0.06 0.89 0.06 0.89 0.315 0.95 0.315 0.95 0.375 0.83 0.375 0.83 0.06 0.3 0.06 0.3 0.405 0.24 0.405 0.24 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.56 0.725 1.035 0.725 1.035 1.055 0.315 1.055 0.315 0.995 0.975 0.995 0.975 0.535 0.68 0.535 0.68 0.515 0.52 0.515 0.52 0.455 0.73 0.455 0.73 0.475 1.035 0.475 1.035 0.665 1.56 0.665 ;
  END
END CLKAND2X4

MACRO CLKAND2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X6 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.437 LAYER Metal1 ;
    ANTENNADIFFAREA 2.001025 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.18803425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 63.82905975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.73 1.37 2.67 1.37 2.67 0.92 2.32 0.92 2.32 1.37 2.26 1.37 2.26 0.92 1.91 0.92 1.91 1.37 1.85 1.37 1.85 0.86 2.46 0.86 2.46 0.585 1.795 0.585 1.795 0.275 1.855 0.275 1.855 0.525 2.205 0.525 2.205 0.275 2.265 0.275 2.265 0.525 2.615 0.525 2.615 0.275 2.675 0.275 2.675 0.585 2.52 0.585 2.52 0.79 2.54 0.79 2.54 0.86 2.73 0.86 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0819 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.893773 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.19 0.895 0.54 0.895 0.54 0.785 0.66 0.785 0.66 0.815 1.07 0.815 1.07 0.785 1.19 0.785 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0819 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.4945055 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.535 0.745 1.475 0.745 1.475 0.685 0.365 0.685 0.365 0.705 0.175 0.705 0.175 0.645 0.235 0.645 0.235 0.625 1.535 0.625 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.28 0.13 1.28 0.13 1.65 0.47 1.65 0.47 1.28 0.53 1.28 0.53 1.65 0.87 1.65 0.87 1.28 0.93 1.28 0.93 1.65 1.2 1.65 1.2 1.28 1.26 1.28 1.26 1.65 1.615 1.65 1.615 1.28 1.675 1.28 1.675 1.65 2.055 1.65 2.055 1.02 2.115 1.02 2.115 1.65 2.465 1.65 2.465 1.02 2.525 1.02 2.525 1.65 2.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 0.06 2.47 0.06 2.47 0.395 2.41 0.395 2.41 0.06 2.06 0.06 2.06 0.395 2 0.395 2 0.06 1.57 0.06 1.57 0.305 1.63 0.305 1.63 0.365 1.51 0.365 1.51 0.06 0.86 0.06 0.86 0.305 0.92 0.305 0.92 0.365 0.8 0.365 0.8 0.06 0.19 0.06 0.19 0.395 0.13 0.395 0.13 0.06 0 0.06 0 -0.06 2.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.22 0.76 1.695 0.76 1.695 1.055 0.205 1.055 0.205 0.995 1.635 0.995 1.635 0.525 0.56 0.525 0.56 0.505 0.49 0.505 0.49 0.445 0.61 0.445 0.61 0.465 1.2 0.465 1.2 0.445 1.32 0.445 1.32 0.465 1.695 0.465 1.695 0.7 2.22 0.7 ;
  END
END CLKAND2X6

MACRO CLKAND2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKAND2X8 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.620575 LAYER Metal1 ;
    ANTENNADIFFAREA 2.422775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.95227375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 52.70270275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.24 1.39 3.18 1.39 3.18 1.005 2.83 1.005 2.83 1.39 2.77 1.39 2.77 1.005 2.42 1.005 2.42 1.39 2.36 1.39 2.36 1.005 2.01 1.005 2.01 1.39 1.95 1.39 1.95 0.945 3.06 0.945 3.06 0.585 1.925 0.585 1.925 0.57 1.865 0.57 1.865 0.51 1.985 0.51 1.985 0.525 2.275 0.525 2.275 0.51 2.395 0.51 2.395 0.525 2.685 0.525 2.685 0.51 2.805 0.51 2.805 0.525 3.08 0.525 3.08 0.51 3.215 0.51 3.215 0.57 3.125 0.57 3.125 0.585 3.12 0.585 3.12 0.79 3.14 0.79 3.14 0.945 3.24 0.945 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0819 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.058608 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.61 0.815 1.365 0.895 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0819 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.5677655 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.605 0.775 1.545 0.775 1.545 0.715 0.235 0.715 0.235 0.625 0.365 0.625 0.365 0.655 1.605 0.655 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 1.77 0 1.77 0 1.65 0.14 1.65 0.14 1.51 0.2 1.51 0.2 1.65 0.54 1.65 0.54 1.51 0.6 1.51 0.6 1.65 0.94 1.65 0.94 1.51 1 1.51 1 1.65 1.35 1.65 1.35 1.51 1.41 1.51 1.41 1.65 1.715 1.65 1.715 1.51 1.775 1.51 1.775 1.65 2.155 1.65 2.155 1.105 2.215 1.105 2.215 1.65 2.565 1.65 2.565 1.105 2.625 1.105 2.625 1.65 2.975 1.65 2.975 1.105 3.035 1.105 3.035 1.65 3.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 0.06 2.98 0.06 2.98 0.425 2.92 0.425 2.92 0.06 2.57 0.06 2.57 0.425 2.51 0.425 2.51 0.06 2.16 0.06 2.16 0.425 2.1 0.425 2.1 0.06 1.65 0.06 1.65 0.335 1.71 0.335 1.71 0.395 1.59 0.395 1.59 0.06 0.94 0.06 0.94 0.335 1 0.335 1 0.395 0.88 0.395 0.88 0.06 0.26 0.06 0.26 0.425 0.2 0.425 0.2 0.06 0 0.06 0 -0.06 3.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.73 0.745 1.765 0.745 1.765 1.055 0.275 1.055 0.275 0.995 1.705 0.995 1.705 0.555 0.64 0.555 0.64 0.535 0.57 0.535 0.57 0.475 0.69 0.475 0.69 0.495 1.28 0.495 1.28 0.475 1.4 0.475 1.4 0.495 1.765 0.495 1.765 0.685 2.73 0.685 ;
  END
END CLKAND2X8

MACRO CLKBUFX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX12 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7804 LAYER Metal1 ;
    ANTENNADIFFAREA 2.4529 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.351 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.07236475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 40.78632475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.98 0.535 0.295 0.535 0.295 0.98 1.98 0.98 1.98 1.45 1.92 1.45 1.92 1.04 1.57 1.04 1.57 1.45 1.51 1.45 1.51 1.04 1.16 1.04 1.16 1.45 1.1 1.45 1.1 1.04 0.75 1.04 0.75 1.45 0.69 1.45 0.69 1.04 0.34 1.04 0.34 1.45 0.26 1.45 0.26 1.04 0.235 1.04 0.235 0.475 0.28 0.475 0.28 0.255 0.34 0.255 0.34 0.475 0.69 0.475 0.69 0.255 0.75 0.255 0.75 0.475 1.1 0.475 1.1 0.255 1.16 0.255 1.16 0.475 1.51 0.475 1.51 0.255 1.57 0.255 1.57 0.475 1.92 0.475 1.92 0.255 1.98 0.255 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.08775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.982906 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.405 0.875 2.34 0.875 2.34 1.23 2.26 1.23 2.26 0.795 2.405 0.795 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.77 0 1.77 0 1.65 0.075 1.65 0.075 0.98 0.135 0.98 0.135 1.65 0.485 1.65 0.485 1.14 0.545 1.14 0.545 1.65 0.895 1.65 0.895 1.14 0.955 1.14 0.955 1.65 1.305 1.65 1.305 1.14 1.365 1.14 1.365 1.65 1.715 1.65 1.715 1.14 1.775 1.14 1.775 1.65 2.125 1.65 2.125 1.33 2.185 1.33 2.185 1.65 2.665 1.65 2.665 1.22 2.725 1.22 2.725 1.65 3 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 0.06 2.725 0.06 2.725 0.425 2.665 0.425 2.665 0.06 2.185 0.06 2.185 0.425 2.125 0.425 2.125 0.06 1.775 0.06 1.775 0.375 1.715 0.375 1.715 0.06 1.365 0.06 1.365 0.375 1.305 0.375 1.305 0.06 0.955 0.06 0.955 0.375 0.895 0.375 0.895 0.06 0.545 0.06 0.545 0.375 0.485 0.375 0.485 0.06 0.135 0.06 0.135 0.565 0.075 0.565 0.075 0.06 0 0.06 0 -0.06 3 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.93 0.695 2.565 0.695 2.565 1.06 2.93 1.06 2.93 1.45 2.87 1.45 2.87 1.12 2.52 1.12 2.52 1.45 2.46 1.45 2.46 1.06 2.505 1.06 2.505 0.695 1.935 0.695 1.935 0.705 1.815 0.705 1.815 0.695 1.54 0.695 1.54 0.705 1.42 0.705 1.42 0.695 1.32 0.695 1.32 0.705 1.2 0.705 1.2 0.695 0.91 0.695 0.91 0.705 0.79 0.705 0.79 0.695 0.69 0.695 0.69 0.705 0.395 0.705 0.395 0.645 0.65 0.645 0.65 0.635 2.46 0.635 2.46 0.445 2.52 0.445 2.52 0.635 2.87 0.635 2.87 0.445 2.93 0.445 ;
  END
END CLKBUFX12

MACRO CLKBUFX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX16 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.378 LAYER Metal1 ;
    ANTENNADIFFAREA 3.1578 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4662 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.100815 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 40.945946 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.825 0.63 2.735 0.63 2.735 0.645 0.29 0.645 0.29 0.905 2.795 0.905 2.795 1.345 2.735 1.345 2.735 0.965 2.385 0.965 2.385 1.345 2.325 1.345 2.325 0.965 1.975 0.965 1.975 1.345 1.915 1.345 1.915 0.965 1.565 0.965 1.565 1.345 1.505 1.345 1.505 0.965 1.155 0.965 1.155 1.345 1.095 1.345 1.095 0.965 0.745 0.965 0.745 1.345 0.685 1.345 0.685 0.965 0.34 0.965 0.34 1.11 0.335 1.11 0.335 1.345 0.26 1.345 0.26 0.965 0.23 0.965 0.23 0.585 0.275 0.585 0.275 0.525 0.335 0.525 0.335 0.585 0.655 0.585 0.655 0.57 0.775 0.57 0.775 0.585 1.065 0.585 1.065 0.57 1.185 0.57 1.185 0.585 1.475 0.585 1.475 0.57 1.595 0.57 1.595 0.585 1.885 0.585 1.885 0.57 2.005 0.57 2.005 0.585 2.295 0.585 2.295 0.57 2.415 0.57 2.415 0.585 2.69 0.585 2.69 0.57 2.825 0.57 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.815 3.76 0.895 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.9 0.13 0.9 0.13 1.65 0.48 1.65 0.48 1.065 0.54 1.065 0.54 1.65 0.89 1.65 0.89 1.065 0.95 1.065 0.95 1.65 1.3 1.65 1.3 1.065 1.36 1.065 1.36 1.65 1.71 1.65 1.71 1.065 1.77 1.065 1.77 1.65 2.12 1.65 2.12 1.065 2.18 1.065 2.18 1.65 2.53 1.65 2.53 1.065 2.59 1.065 2.59 1.65 2.94 1.65 2.94 0.955 3 0.955 3 1.65 3.35 1.65 3.35 1.225 3.41 1.225 3.41 1.65 3.86 1.65 3.86 0.955 3.92 0.955 3.92 1.65 4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.82 0.06 3.82 0.52 3.76 0.52 3.76 0.06 3.41 0.06 3.41 0.52 3.35 0.52 3.35 0.06 3 0.06 3 0.52 2.94 0.52 2.94 0.06 2.59 0.06 2.59 0.485 2.53 0.485 2.53 0.06 2.18 0.06 2.18 0.485 2.12 0.485 2.12 0.06 1.77 0.06 1.77 0.485 1.71 0.485 1.71 0.06 1.36 0.06 1.36 0.485 1.3 0.485 1.3 0.06 0.95 0.06 0.95 0.485 0.89 0.485 0.89 0.06 0.54 0.06 0.54 0.485 0.48 0.485 0.48 0.06 0.13 0.06 0.13 0.485 0.07 0.485 0.07 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.615 0.68 3.16 0.68 3.16 0.995 3.615 0.995 3.615 1.345 3.555 1.345 3.555 1.055 3.205 1.055 3.205 1.345 3.145 1.345 3.145 1.055 3.1 1.055 3.1 0.805 0.39 0.805 0.39 0.745 3.1 0.745 3.1 0.62 3.145 0.62 3.145 0.54 3.205 0.54 3.205 0.62 3.555 0.62 3.555 0.54 3.615 0.54 ;
  END
END CLKBUFX16

MACRO CLKBUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX2 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4428 LAYER Metal1 ;
    ANTENNADIFFAREA 0.6098 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.56923075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 63.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.41 0.615 0.365 0.615 0.365 0.865 0.41 0.865 0.41 1.32 0.35 1.32 0.35 0.925 0.305 0.925 0.305 0.73 0.26 0.73 0.26 0.6 0.305 0.6 0.305 0.555 0.35 0.555 0.35 0.495 0.41 0.495 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.765 1.085 0.51 1.085 0.51 1.005 0.685 1.005 0.685 0.76 0.765 0.76 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.145 1.65 0.145 0.93 0.205 0.93 0.205 1.65 0.555 1.65 0.555 1.185 0.615 1.185 0.615 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.615 0.06 0.615 0.5 0.555 0.5 0.555 0.06 0.205 0.06 0.205 0.5 0.145 0.5 0.145 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.925 1.21 0.865 1.21 0.865 0.66 0.585 0.66 0.585 0.77 0.465 0.77 0.465 0.71 0.525 0.71 0.525 0.6 0.865 0.6 0.865 0.405 0.925 0.405 ;
  END
END CLKBUFX2

MACRO CLKBUFX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX20 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.97005 LAYER Metal1 ;
    ANTENNADIFFAREA 3.839 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.0770085 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 41.076923 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.41 0.655 0.14 0.655 0.14 0.915 3.41 0.915 3.41 1.36 3.35 1.36 3.35 0.975 3 0.975 3 1.36 2.94 1.36 2.94 0.975 2.59 0.975 2.59 1.36 2.53 1.36 2.53 0.975 2.18 0.975 2.18 1.36 2.12 1.36 2.12 0.975 1.77 0.975 1.77 1.36 1.71 1.36 1.71 0.975 1.36 0.975 1.36 1.36 1.3 1.36 1.3 0.975 0.95 0.975 0.95 1.36 0.89 1.36 0.89 0.975 0.54 0.975 0.54 1.36 0.48 1.36 0.48 0.975 0.13 0.975 0.13 1.36 0.06 1.36 0.06 0.355 0.13 0.355 0.13 0.595 0.48 0.595 0.48 0.355 0.54 0.355 0.54 0.595 0.89 0.595 0.89 0.355 0.95 0.355 0.95 0.595 1.3 0.595 1.3 0.355 1.36 0.355 1.36 0.595 1.71 0.595 1.71 0.355 1.77 0.355 1.77 0.595 2.12 0.595 2.12 0.355 2.18 0.355 2.18 0.595 2.53 0.595 2.53 0.355 2.59 0.355 2.59 0.595 2.94 0.595 2.94 0.355 3 0.355 3 0.595 3.35 0.595 3.35 0.355 3.41 0.355 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.14625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.1897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.875 0.815 4.375 0.895 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.075 0.335 1.075 0.335 1.65 0.685 1.65 0.685 1.075 0.745 1.075 0.745 1.65 1.095 1.65 1.095 1.075 1.155 1.075 1.155 1.65 1.505 1.65 1.505 1.075 1.565 1.075 1.565 1.65 1.915 1.65 1.915 1.075 1.975 1.075 1.975 1.65 2.325 1.65 2.325 1.075 2.385 1.075 2.385 1.65 2.735 1.65 2.735 1.075 2.795 1.075 2.795 1.65 3.145 1.65 3.145 1.075 3.205 1.075 3.205 1.65 3.555 1.65 3.555 0.97 3.615 0.97 3.615 1.65 3.965 1.65 3.965 1.24 4.025 1.24 4.025 1.65 4.375 1.65 4.375 1.24 4.435 1.24 4.435 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 4.435 0.06 4.435 0.52 4.375 0.52 4.375 0.06 4.025 0.06 4.025 0.52 3.965 0.52 3.965 0.06 3.615 0.06 3.615 0.52 3.555 0.52 3.555 0.06 3.205 0.06 3.205 0.475 3.145 0.475 3.145 0.06 2.795 0.06 2.795 0.475 2.735 0.475 2.735 0.06 2.385 0.06 2.385 0.475 2.325 0.475 2.325 0.06 1.975 0.06 1.975 0.475 1.915 0.475 1.915 0.06 1.565 0.06 1.565 0.475 1.505 0.475 1.505 0.06 1.155 0.06 1.155 0.475 1.095 0.475 1.095 0.06 0.745 0.06 0.745 0.475 0.685 0.475 0.685 0.06 0.335 0.06 0.335 0.475 0.275 0.475 0.275 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.64 0.68 3.775 0.68 3.775 0.995 4.64 0.995 4.64 1.36 4.58 1.36 4.58 1.055 4.23 1.055 4.23 1.36 4.17 1.36 4.17 1.055 3.82 1.055 3.82 1.36 3.76 1.36 3.76 1.055 3.715 1.055 3.715 0.815 0.31 0.815 0.31 0.755 3.715 0.755 3.715 0.62 3.76 0.62 3.76 0.54 3.82 0.54 3.82 0.62 4.17 0.62 4.17 0.54 4.23 0.54 4.23 0.62 4.58 0.62 4.58 0.54 4.64 0.54 ;
  END
END CLKBUFX20

MACRO CLKBUFX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX3 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6117 LAYER Metal1 ;
    ANTENNADIFFAREA 0.79045 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.08775 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.97094025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 55.4188035 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.685 1.44 0.625 1.44 0.625 1.11 0.275 1.11 0.275 1.44 0.215 1.44 0.215 1.05 0.26 1.05 0.26 0.62 0.175 0.62 0.175 0.48 0.235 0.48 0.235 0.56 0.54 0.56 0.54 0.405 0.585 0.405 0.585 0.345 0.645 0.345 0.645 0.465 0.6 0.465 0.6 0.62 0.32 0.62 0.32 0.98 0.34 0.98 0.34 1.05 0.685 1.05 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.72 0.94 1.22 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.42 1.65 0.42 1.21 0.48 1.21 0.48 1.65 0.83 1.65 0.83 1.32 0.89 1.32 0.89 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.85 0.06 0.85 0.46 0.79 0.46 0.79 0.06 0.44 0.06 0.44 0.46 0.38 0.46 0.38 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.1 1.44 1.04 1.44 1.04 0.62 0.76 0.62 0.76 0.77 0.7 0.77 0.7 0.56 1.02 0.56 1.02 0.48 1.1 0.48 ;
  END
END CLKBUFX3

MACRO CLKBUFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX4 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.795775 LAYER Metal1 ;
    ANTENNADIFFAREA 0.94375 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.80149575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 54.4102565 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 0.48 0.305 0.48 0.305 0.905 0.76 0.905 0.76 1.37 0.7 1.37 0.7 0.965 0.335 0.965 0.335 1.37 0.275 1.37 0.275 0.965 0.23 0.965 0.23 0.84 0.225 0.84 0.225 0.76 0.23 0.76 0.23 0.42 0.275 0.42 0.275 0.23 0.335 0.23 0.335 0.42 0.7 0.42 0.7 0.23 0.76 0.23 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.051282 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.03 0.86 0.94 0.86 0.94 0.965 0.86 0.965 0.86 0.74 1.03 0.74 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.98 0.13 0.98 0.13 1.65 0.48 1.65 0.48 1.095 0.54 1.095 0.54 1.65 0.905 1.65 0.905 1.095 0.965 1.095 0.965 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 0.965 0.06 0.965 0.48 0.905 0.48 0.905 0.06 0.54 0.06 0.54 0.36 0.48 0.36 0.48 0.06 0.13 0.06 0.13 0.48 0.07 0.48 0.07 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.175 1.37 1.11 1.37 1.11 0.64 0.39 0.64 0.39 0.58 1.11 0.58 1.11 0.23 1.175 0.23 ;
  END
END CLKBUFX4

MACRO CLKBUFX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX6 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.565 0.06 1.565 0.47 1.505 0.47 1.505 0.06 1.155 0.06 1.155 0.47 1.095 0.47 1.095 0.06 0.745 0.06 0.745 0.47 0.685 0.47 0.685 0.06 0.335 0.06 0.335 0.47 0.275 0.47 0.275 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.075 0.335 1.075 0.335 1.65 0.685 1.65 0.685 1.075 0.745 1.075 0.745 1.65 1.095 1.65 1.095 0.915 1.155 0.915 1.155 1.65 1.505 1.65 1.505 1.17 1.565 1.17 1.565 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.57 1.54 1.07 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02695 LAYER Metal1 ;
    ANTENNADIFFAREA 1.3524 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.851567 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 46.82051275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.95 0.655 0.13 0.655 0.13 0.79 0.14 0.79 0.14 0.915 0.95 0.915 0.95 1.37 0.89 1.37 0.89 0.975 0.54 0.975 0.54 1.37 0.48 1.37 0.48 0.975 0.13 0.975 0.13 1.37 0.06 1.37 0.06 0.35 0.13 0.35 0.13 0.595 0.48 0.595 0.48 0.35 0.54 0.35 0.54 0.595 0.89 0.595 0.89 0.35 0.95 0.35 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      POLYGON 1.36 1.29 1.3 1.29 1.3 0.815 0.32 0.815 0.32 0.755 1.3 0.755 1.3 0.49 1.36 0.49 ;
  END
END CLKBUFX6

MACRO CLKBUFX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKBUFX8 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3434 LAYER Metal1 ;
    ANTENNADIFFAREA 1.65 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.76319175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 46.988417 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.515 0.705 0.305 0.705 0.305 0.93 1.515 0.93 1.515 1.375 1.455 1.375 1.455 0.99 1.105 0.99 1.105 1.375 1.045 1.375 1.045 0.99 0.695 0.99 0.695 1.375 0.635 1.375 0.635 0.99 0.285 0.99 0.285 1.375 0.225 1.375 0.225 0.345 0.285 0.345 0.285 0.645 0.635 0.645 0.635 0.345 0.695 0.345 0.695 0.645 1.045 0.645 1.045 0.345 1.105 0.345 1.105 0.645 1.455 0.645 1.455 0.345 1.515 0.345 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.74358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2 0.68 2.13 0.89 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.43 1.65 0.43 1.09 0.49 1.09 0.49 1.65 0.84 1.65 0.84 1.09 0.9 1.09 0.9 1.65 1.25 1.65 1.25 1.09 1.31 1.09 1.31 1.65 1.66 1.65 1.66 0.93 1.72 0.93 1.72 1.65 2.07 1.65 2.07 1.06 2.13 1.06 2.13 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 2.13 0.06 2.13 0.62 2.07 0.62 2.07 0.06 1.72 0.06 1.72 0.64 1.66 0.64 1.66 0.06 1.31 0.06 1.31 0.585 1.25 0.585 1.25 0.06 0.9 0.06 0.9 0.585 0.84 0.585 0.84 0.06 0.49 0.06 0.49 0.585 0.43 0.585 0.43 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.925 1.32 1.865 1.32 1.865 0.825 0.54 0.825 0.54 0.765 1.865 0.765 1.865 0.38 1.925 0.38 ;
  END
END CLKBUFX8

MACRO CLKINVX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX1 0 0 ;
  SIZE 0.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2202 LAYER Metal1 ;
    ANTENNADIFFAREA 0.3144 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.335 1.14 0.275 1.14 0.275 0.73 0.255 0.73 0.255 0.6 0.275 0.6 0.275 0.51 0.335 0.51 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.3846155 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.055 0.67 0.19 0.865 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.93 0.13 0.93 0.13 1.65 0.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 0.06 0.13 0.06 0.13 0.61 0.07 0.61 0.07 0.06 0 0.06 0 -0.06 0.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END CLKINVX1

MACRO CLKINVX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX12 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3369 LAYER Metal1 ;
    ANTENNADIFFAREA 2.0307 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.165 0.96 2.14 0.96 2.14 1.37 2.06 1.37 2.06 0.96 1.62 0.96 1.62 1.37 1.56 1.37 1.56 0.96 1.21 0.96 1.21 1.37 1.15 1.37 1.15 0.96 0.8 0.96 0.8 1.37 0.74 1.37 0.74 0.96 0.335 0.96 0.335 1.37 0.275 1.37 0.275 0.9 2.105 0.9 2.105 0.525 0.33 0.525 0.33 0.23 0.39 0.23 0.39 0.465 0.74 0.465 0.74 0.23 0.8 0.23 0.8 0.465 1.15 0.465 1.15 0.23 1.21 0.23 1.21 0.465 1.56 0.465 1.56 0.23 1.62 0.23 1.62 0.465 1.99 0.465 1.99 0.23 2.05 0.23 2.05 0.465 2.165 0.465 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.351 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4615385 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.005 0.685 0.565 0.685 0.565 0.705 0.435 0.705 0.435 0.685 0.375 0.685 0.375 0.625 2.005 0.625 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.9 0.13 0.9 0.13 1.65 0.48 1.65 0.48 1.25 0.54 1.25 0.54 1.65 0.945 1.65 0.945 1.25 1.005 1.25 1.005 1.65 1.355 1.65 1.355 1.25 1.415 1.25 1.415 1.65 1.765 1.65 1.765 1.25 1.825 1.25 1.825 1.65 2.265 1.65 2.265 0.9 2.325 0.9 2.325 1.65 2.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 0.06 2.325 0.06 2.325 0.54 2.265 0.54 2.265 0.06 1.845 0.06 1.845 0.35 1.785 0.35 1.785 0.06 1.415 0.06 1.415 0.35 1.355 0.35 1.355 0.06 1.005 0.06 1.005 0.35 0.945 0.35 0.945 0.06 0.595 0.06 0.595 0.35 0.535 0.35 0.535 0.06 0.13 0.06 0.13 0.54 0.07 0.54 0.07 0.06 0 0.06 0 -0.06 2.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END CLKINVX12

MACRO CLKINVX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX16 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.215 LAYER Metal1 ;
    ANTENNADIFFAREA 2.5144 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.97 0.99 2.94 0.99 2.94 1.11 2.925 1.11 2.925 1.345 2.865 1.345 2.865 1.11 2.86 1.11 2.86 0.99 2.515 0.99 2.515 1.345 2.455 1.345 2.455 0.99 2.105 0.99 2.105 1.345 2.045 1.345 2.045 0.99 1.695 0.99 1.695 1.345 1.635 1.345 1.635 1.055 1.285 1.055 1.285 1.345 1.225 1.345 1.225 1.055 0.895 1.055 0.895 1.345 0.815 1.345 0.815 1.055 0.465 1.055 0.465 1.345 0.405 1.345 0.405 0.995 1.635 0.995 1.635 0.93 2.91 0.93 2.91 0.645 0.45 0.645 0.45 0.63 0.375 0.63 0.375 0.57 0.495 0.57 0.495 0.585 0.785 0.585 0.785 0.57 0.905 0.57 0.905 0.585 1.195 0.585 1.195 0.57 1.315 0.57 1.315 0.585 1.605 0.585 1.605 0.57 1.725 0.57 1.725 0.585 2.015 0.585 2.015 0.57 2.135 0.57 2.135 0.585 2.425 0.585 2.425 0.57 2.545 0.57 2.545 0.585 2.865 0.585 2.865 0.525 2.925 0.525 2.925 0.585 2.97 0.585 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4662 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.5572715 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.81 0.83 0.765 0.83 0.765 0.895 0.635 0.895 0.635 0.83 0.515 0.83 0.515 0.77 2.81 0.77 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 1.77 0 1.77 0 1.65 0.2 1.65 0.2 0.9 0.26 0.9 0.26 1.65 0.61 1.65 0.61 1.225 0.67 1.225 0.67 1.65 1.02 1.65 1.02 1.225 1.08 1.225 1.08 1.65 1.43 1.65 1.43 1.225 1.49 1.225 1.49 1.65 1.84 1.65 1.84 1.225 1.9 1.225 1.9 1.65 2.25 1.65 2.25 1.225 2.31 1.225 2.31 1.65 2.66 1.65 2.66 1.225 2.72 1.225 2.72 1.65 3.07 1.65 3.07 0.9 3.13 0.9 3.13 1.65 3.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 0.06 3.13 0.06 3.13 0.485 3.07 0.485 3.07 0.06 2.72 0.06 2.72 0.485 2.66 0.485 2.66 0.06 2.31 0.06 2.31 0.485 2.25 0.485 2.25 0.06 1.9 0.06 1.9 0.485 1.84 0.485 1.84 0.06 1.49 0.06 1.49 0.485 1.43 0.485 1.43 0.06 1.08 0.06 1.08 0.485 1.02 0.485 1.02 0.06 0.67 0.06 0.67 0.485 0.61 0.485 0.61 0.06 0.26 0.06 0.26 0.485 0.2 0.485 0.2 0.06 0 0.06 0 -0.06 3.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END CLKINVX16

MACRO CLKINVX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX2 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3348 LAYER Metal1 ;
    ANTENNADIFFAREA 0.478 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.52 0.54 1.29 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.36 0.8 0.28 0.8 0.28 0.76 0.06 0.76 0.06 0.6 0.14 0.6 0.14 0.68 0.28 0.68 0.28 0.6 0.36 0.6 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.77 0 1.77 0 1.65 0.255 1.65 0.255 0.9 0.315 0.9 0.315 1.65 0.665 1.65 0.665 0.9 0.725 0.9 0.725 1.65 0.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 0.06 0.725 0.06 0.725 0.5 0.665 0.5 0.665 0.06 0.315 0.06 0.315 0.5 0.255 0.5 0.255 0.06 0 0.06 0 -0.06 0.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END CLKINVX2

MACRO CLKINVX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX20 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1593 LAYER Metal1 ;
    ANTENNADIFFAREA 3.122275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.7 1.36 3.64 1.36 3.64 0.98 3.205 0.98 3.205 1.36 3.145 1.36 3.145 0.98 2.795 0.98 2.795 1.36 2.735 1.36 2.735 0.98 2.385 0.98 2.385 1.36 2.325 1.36 2.325 0.98 1.975 0.98 1.975 1.36 1.915 1.36 1.915 0.98 1.565 0.98 1.565 1.36 1.505 1.36 1.505 0.98 1.155 0.98 1.155 1.36 1.095 1.36 1.095 1.14 0.745 1.14 0.745 1.36 0.685 1.36 0.685 1.14 0.335 1.14 0.335 1.36 0.275 1.36 0.275 0.92 0.335 0.92 0.335 1.08 0.685 1.08 0.685 0.92 0.745 0.92 0.745 1.08 1.095 1.08 1.095 0.92 3.3 0.92 3.3 0.66 0.275 0.66 0.275 0.355 0.335 0.355 0.335 0.6 0.685 0.6 0.685 0.355 0.745 0.355 0.745 0.6 1.095 0.6 1.095 0.355 1.155 0.355 1.155 0.6 1.505 0.6 1.505 0.355 1.565 0.355 1.565 0.6 1.915 0.6 1.915 0.355 1.975 0.355 1.975 0.6 2.325 0.6 2.325 0.355 2.385 0.355 2.385 0.6 2.735 0.6 2.735 0.355 2.795 0.355 2.795 0.6 3.145 0.6 3.145 0.355 3.205 0.355 3.205 0.6 3.555 0.6 3.555 0.355 3.615 0.355 3.615 0.66 3.36 0.66 3.36 0.92 3.46 0.92 3.46 0.79 3.54 0.79 3.54 0.92 3.64 0.92 3.64 0.905 3.7 0.905 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.497436 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.105 0.82 0.565 0.82 0.565 0.895 0.435 0.895 0.435 0.82 0.32 0.82 0.32 0.76 3.105 0.76 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.9 0.13 0.9 0.13 1.65 0.48 1.65 0.48 1.24 0.54 1.24 0.54 1.65 0.89 1.65 0.89 1.24 0.95 1.24 0.95 1.65 1.3 1.65 1.3 1.24 1.36 1.24 1.36 1.65 1.71 1.65 1.71 1.24 1.77 1.24 1.77 1.65 2.12 1.65 2.12 1.24 2.18 1.24 2.18 1.65 2.53 1.65 2.53 1.24 2.59 1.24 2.59 1.65 2.94 1.65 2.94 1.24 3 1.24 3 1.65 3.35 1.65 3.35 1.24 3.41 1.24 3.41 1.65 3.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 0.06 3.41 0.06 3.41 0.475 3.35 0.475 3.35 0.06 3 0.06 3 0.475 2.94 0.475 2.94 0.06 2.59 0.06 2.59 0.475 2.53 0.475 2.53 0.06 2.18 0.06 2.18 0.475 2.12 0.475 2.12 0.06 1.77 0.06 1.77 0.475 1.71 0.475 1.71 0.06 1.36 0.06 1.36 0.475 1.3 0.475 1.3 0.06 0.95 0.06 0.95 0.475 0.89 0.475 0.89 0.06 0.54 0.06 0.54 0.475 0.48 0.475 0.48 0.06 0.13 0.06 0.13 0.66 0.07 0.66 0.07 0.06 0 0.06 0 -0.06 3.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END CLKINVX20

MACRO CLKINVX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX3 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3669 LAYER Metal1 ;
    ANTENNADIFFAREA 0.63 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.885 0.68 0.54 0.68 0.54 0.9 0.885 0.9 0.885 1.29 0.825 1.29 0.825 0.96 0.475 0.96 0.475 1.29 0.415 1.29 0.415 0.9 0.46 0.9 0.46 0.68 0.415 0.68 0.415 0.54 0.475 0.54 0.475 0.62 0.825 0.62 0.825 0.54 0.885 0.54 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.08775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.982906 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.315 0.945 0.06 0.945 0.06 0.725 0.235 0.725 0.235 0.62 0.315 0.62 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.21 1.65 0.21 1.045 0.27 1.045 0.27 1.65 0.62 1.65 0.62 1.06 0.68 1.06 0.68 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.68 0.06 0.68 0.52 0.62 0.52 0.62 0.06 0.27 0.06 0.27 0.52 0.21 0.52 0.21 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END CLKINVX3

MACRO CLKINVX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX4 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.422725 LAYER Metal1 ;
    ANTENNADIFFAREA 0.763375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.815 1.11 0.745 1.11 0.745 1.335 0.685 1.335 0.685 1.015 0.335 1.015 0.335 1.335 0.275 1.335 0.275 0.955 0.735 0.955 0.735 0.755 0.275 0.755 0.275 0.415 0.335 0.415 0.335 0.695 0.685 0.695 0.685 0.415 0.745 0.415 0.745 0.695 0.795 0.695 0.795 0.98 0.815 0.98 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.32051275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.2 0.815 0.635 0.895 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.945 0.13 0.945 0.13 1.65 0.48 1.65 0.48 1.095 0.54 1.095 0.54 1.65 0.815 1.65 0.815 1.51 0.94 1.51 0.94 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.94 0.06 0.94 0.225 0.815 0.225 0.815 0.06 0.54 0.06 0.54 0.635 0.48 0.635 0.48 0.06 0.13 0.06 0.13 0.635 0.07 0.635 0.07 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END CLKINVX4

MACRO CLKINVX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX6 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7396 LAYER Metal1 ;
    ANTENNADIFFAREA 1.0614 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.165 0.525 0.92 0.525 0.92 0.79 0.94 0.79 0.94 0.9 1.165 0.9 1.165 1.37 1.105 1.37 1.105 0.96 0.755 0.96 0.755 1.37 0.695 1.37 0.695 1.15 0.335 1.15 0.335 1.37 0.275 1.37 0.275 0.9 0.335 0.9 0.335 1.09 0.695 1.09 0.695 0.9 0.86 0.9 0.86 0.525 0.285 0.525 0.285 0.245 0.345 0.245 0.345 0.465 0.695 0.465 0.695 0.245 0.755 0.245 0.755 0.465 1.105 0.465 1.105 0.245 1.165 0.245 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 0.991453 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.625 0.73 0.705 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.9 0.13 0.9 0.13 1.65 0.48 1.65 0.48 1.25 0.54 1.25 0.54 1.65 0.9 1.65 0.9 1.25 0.96 1.25 0.96 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 0.96 0.06 0.96 0.365 0.9 0.365 0.9 0.06 0.55 0.06 0.55 0.365 0.49 0.365 0.49 0.06 0.13 0.06 0.13 0.555 0.07 0.555 0.07 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END CLKINVX6

MACRO CLKINVX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKINVX8 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6555 LAYER Metal1 ;
    ANTENNADIFFAREA 1.3496 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.645 0.63 1.57 0.63 1.57 0.645 1.34 0.645 1.34 0.73 1.32 0.73 1.32 0.96 1.615 0.96 1.615 1.345 1.555 1.345 1.555 1.02 1.205 1.02 1.205 1.345 1.145 1.345 1.145 1.055 0.795 1.055 0.795 1.345 0.735 1.345 0.735 1.055 0.385 1.055 0.385 1.345 0.325 1.345 0.325 0.995 1.135 0.995 1.135 0.96 1.26 0.96 1.26 0.645 0.37 0.645 0.37 0.63 0.295 0.63 0.295 0.57 0.415 0.57 0.415 0.585 0.705 0.585 0.705 0.57 0.825 0.57 0.825 0.585 1.145 0.585 1.145 0.525 1.205 0.525 1.205 0.585 1.525 0.585 1.525 0.57 1.645 0.57 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.010296 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.095 0.85 0.565 0.85 0.565 0.895 0.435 0.895 0.435 0.77 1.095 0.77 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.12 1.65 0.12 0.9 0.18 0.9 0.18 1.65 0.53 1.65 0.53 1.225 0.59 1.225 0.59 1.65 0.94 1.65 0.94 1.225 1 1.225 1 1.65 1.35 1.65 1.35 1.225 1.41 1.225 1.41 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.41 0.06 1.41 0.485 1.35 0.485 1.35 0.06 1 0.06 1 0.485 0.94 0.485 0.94 0.06 0.59 0.06 0.59 0.485 0.53 0.485 0.53 0.06 0.18 0.06 0.18 0.485 0.12 0.485 0.12 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END CLKINVX8

MACRO CLKMX2X12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X12 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.06805 LAYER Metal1 ;
    ANTENNADIFFAREA 2.7787 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.374175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.52695925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 43.53577875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.335 1.48 3.275 1.48 3.275 0.98 3.23 0.98 3.23 0.85 2.925 0.85 2.925 1.48 2.865 1.48 2.865 0.85 2.515 0.85 2.515 1.48 2.455 1.48 2.455 0.85 2.105 0.85 2.105 1.48 2.045 1.48 2.045 0.85 1.74 0.85 1.74 0.92 1.695 0.92 1.695 1.48 1.635 1.48 1.635 0.535 1.54 0.535 1.54 0.415 1.6 0.415 1.6 0.475 1.695 0.475 1.695 0.79 2 0.79 2 0.3 2.06 0.3 2.06 0.79 2.41 0.79 2.41 0.3 2.47 0.3 2.47 0.79 2.82 0.79 2.82 0.3 2.88 0.3 2.88 0.79 3.23 0.79 3.23 0.3 3.29 0.3 3.29 0.92 3.335 0.92 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 1.11 1.305 1.11 1.305 1.26 1.225 1.26 1.225 0.99 1.26 0.99 1.26 0.795 1.34 0.795 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.472492 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.68 0.56 1.08 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.052425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.8941345 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.805 1.115 0.74 1.115 0.74 1.26 0.26 1.26 0.26 0.92 0.34 0.92 0.34 1.18 0.66 1.18 0.66 1.035 0.805 1.035 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 1.77 0 1.77 0 1.65 0.425 1.65 0.425 1.36 0.485 1.36 0.485 1.65 1.43 1.65 1.43 1.36 1.49 1.36 1.49 1.65 1.84 1.65 1.84 1.01 1.9 1.01 1.9 1.65 2.25 1.65 2.25 1.01 2.31 1.01 2.31 1.65 2.66 1.65 2.66 1.01 2.72 1.01 2.72 1.65 3.07 1.65 3.07 1.01 3.13 1.01 3.13 1.65 3.48 1.65 3.48 1.01 3.54 1.01 3.54 1.65 3.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 0.06 3.495 0.06 3.495 0.61 3.435 0.61 3.435 0.06 3.085 0.06 3.085 0.61 3.025 0.61 3.025 0.06 2.675 0.06 2.675 0.61 2.615 0.61 2.615 0.06 2.265 0.06 2.265 0.61 2.205 0.61 2.205 0.06 1.855 0.06 1.855 0.61 1.795 0.61 1.795 0.06 1.36 0.06 1.36 0.42 1.3 0.42 1.3 0.06 0.485 0.06 0.485 0.42 0.425 0.42 0.425 0.06 0 0.06 0 -0.06 3.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.535 0.795 1.475 0.795 1.475 0.695 1.125 0.695 1.125 1.275 0.9 1.275 0.9 1.335 0.84 1.335 0.84 1.215 1.065 1.215 1.065 0.42 0.735 0.42 0.735 0.3 0.795 0.3 0.795 0.36 1.125 0.36 1.125 0.635 1.535 0.635 ;
      POLYGON 0.965 1.115 0.905 1.115 0.905 0.855 0.72 0.855 0.72 0.665 0.66 0.665 0.66 0.58 0.16 0.58 0.16 1.36 0.28 1.36 0.28 1.48 0.22 1.48 0.22 1.42 0.1 1.42 0.1 0.52 0.22 0.52 0.22 0.44 0.28 0.44 0.28 0.52 0.78 0.52 0.78 0.795 0.965 0.795 ;
  END
END CLKMX2X12

MACRO CLKMX2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8535 LAYER Metal1 ;
    ANTENNADIFFAREA 1.0052 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0747 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.42570275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 91.88755025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 0.73 1.66 0.73 1.66 0.66 1.56 0.66 1.56 1.105 1.525 1.105 1.525 1.435 1.465 1.435 1.465 1.045 1.5 1.045 1.5 0.485 1.465 0.485 1.465 0.365 1.525 0.365 1.525 0.425 1.56 0.425 1.56 0.6 1.74 0.6 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.895 1.3 0.895 1.3 1.215 1.22 1.215 1.22 0.815 1.4 0.815 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.035 0.44 1.035 0.44 0.955 0.46 0.955 0.46 0.635 0.54 0.635 0.54 0.955 0.62 0.955 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.074074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.215 0.26 1.215 0.26 0.98 0.34 0.98 0.34 1.135 0.72 1.135 0.72 0.93 0.8 0.93 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.41 1.65 0.41 1.315 0.47 1.315 0.47 1.65 1.26 1.65 1.26 1.315 1.32 1.315 1.32 1.65 1.67 1.65 1.67 1.045 1.73 1.045 1.73 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.73 0.06 1.73 0.375 1.67 0.375 1.67 0.06 1.32 0.06 1.32 0.375 1.26 0.375 1.26 0.06 0.47 0.06 0.47 0.375 0.41 0.375 0.41 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.4 0.645 1.12 0.645 1.12 1.335 0.89 1.335 0.89 1.275 1.06 1.275 1.06 0.375 0.735 0.375 0.735 0.255 0.795 0.255 0.795 0.315 1.12 0.315 1.12 0.585 1.4 0.585 ;
      POLYGON 0.96 1.155 0.9 1.155 0.9 0.805 0.64 0.805 0.64 0.535 0.16 0.535 0.16 1.315 0.265 1.315 0.265 1.435 0.205 1.435 0.205 1.375 0.1 1.375 0.1 0.475 0.205 0.475 0.205 0.28 0.265 0.28 0.265 0.475 0.76 0.475 0.76 0.745 0.96 0.745 ;
  END
END CLKMX2X2

MACRO CLKMX2X3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X3 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.10925 LAYER Metal1 ;
    ANTENNADIFFAREA 1.603975 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.48076925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 71.897436 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.23 0.58 1.865 0.58 1.865 0.79 1.94 0.79 1.94 0.86 2.23 0.86 2.23 1.365 2.17 1.365 2.17 0.92 1.865 0.92 1.865 1.055 1.82 1.055 1.82 1.365 1.76 1.365 1.76 0.995 1.805 0.995 1.805 0.53 1.73 0.53 1.73 0.47 1.865 0.47 1.865 0.52 2.17 0.52 2.17 0.44 2.23 0.44 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.705 0.895 1.515 0.895 1.515 1.1 1.435 1.1 1.435 0.79 1.515 0.79 1.515 0.815 1.705 0.815 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.795 1.015 0.635 1.015 0.635 0.87 0.44 0.87 0.44 0.79 0.795 0.79 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.339934 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.015 0.9 0.955 0.9 0.955 1.175 0.28 1.175 0.28 0.92 0.26 0.92 0.26 0.79 0.34 0.79 0.34 1.115 0.895 1.115 0.895 0.84 1.015 0.84 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 1.77 0 1.77 0 1.65 0.65 1.65 0.65 1.275 0.77 1.275 0.77 1.335 0.71 1.335 0.71 1.65 1.475 1.65 1.475 1.2 1.535 1.2 1.535 1.65 1.965 1.65 1.965 1.02 2.025 1.02 2.025 1.65 2.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 0.06 2.025 0.06 2.025 0.42 1.965 0.42 1.965 0.06 1.535 0.06 1.535 0.42 1.475 0.42 1.475 0.06 0.415 0.06 0.415 0.53 0.355 0.53 0.355 0.06 0 0.06 0 -0.06 2.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.705 0.69 1.335 0.69 1.335 1.06 1.125 1.06 1.125 1.365 1.065 1.365 1.065 1 1.275 1 1.275 0.53 0.875 0.53 0.875 0.47 1.335 0.47 1.335 0.63 1.705 0.63 ;
      POLYGON 1.175 0.9 1.115 0.9 1.115 0.69 0.16 0.69 0.16 1.02 0.18 1.02 0.18 1.14 0.12 1.14 0.12 1.08 0.1 1.08 0.1 0.63 0.15 0.63 0.15 0.435 0.21 0.435 0.21 0.63 1.175 0.63 ;
  END
END CLKMX2X3

MACRO CLKMX2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X4 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1918 LAYER Metal1 ;
    ANTENNADIFFAREA 1.505125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.140175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.50222925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 64.05564475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.995 0.53 1.63 0.53 1.63 0.98 1.74 0.98 1.74 1.05 1.995 1.05 1.995 1.48 1.935 1.48 1.935 1.11 1.585 1.11 1.585 1.48 1.525 1.48 1.525 1.05 1.57 1.05 1.57 0.48 1.495 0.48 1.495 0.42 1.63 0.42 1.63 0.47 1.935 0.47 1.935 0.39 1.995 0.39 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.47 0.895 1.315 0.895 1.315 1.105 1.18 1.105 1.18 0.95 1.235 0.95 1.235 0.815 1.47 0.815 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.63 0.54 1.13 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.039375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.60952375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 0.97 0.7 0.97 0.7 1.29 0.26 1.29 0.26 0.98 0.34 0.98 0.34 1.23 0.64 1.23 0.64 0.91 0.76 0.91 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 1.77 0 1.77 0 1.65 0.395 1.65 0.395 1.39 0.515 1.39 0.515 1.65 1.24 1.65 1.24 1.205 1.3 1.205 1.3 1.65 1.73 1.65 1.73 1.21 1.79 1.21 1.79 1.65 2.14 1.65 2.14 1.09 2.2 1.09 2.2 1.65 2.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 0.06 2.2 0.06 2.2 0.37 2.14 0.37 2.14 0.06 1.79 0.06 1.79 0.37 1.73 0.37 1.73 0.06 1.27 0.06 1.27 0.28 1.33 0.28 1.33 0.34 1.21 0.34 1.21 0.06 0.5 0.06 0.5 0.37 0.44 0.37 0.44 0.06 0 0.06 0 -0.06 2.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.47 0.715 1.08 0.715 1.08 1.265 0.87 1.265 0.87 1.325 0.81 1.325 0.81 1.205 1.02 1.205 1.02 0.37 0.87 0.37 0.87 0.25 0.93 0.25 0.93 0.31 1.08 0.31 1.08 0.655 1.47 0.655 ;
      POLYGON 0.92 1.105 0.86 1.105 0.86 0.66 0.8 0.66 0.8 0.53 0.16 0.53 0.16 1.39 0.295 1.39 0.295 1.45 0.1 1.45 0.1 0.47 0.205 0.47 0.205 0.335 0.265 0.335 0.265 0.47 0.92 0.47 ;
  END
END CLKMX2X4

MACRO CLKMX2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X6 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3599 LAYER Metal1 ;
    ANTENNADIFFAREA 1.815075 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.198675 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.844847 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 53.7561345 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.515 1.395 2.455 1.395 2.455 0.985 2.41 0.985 2.41 0.66 2.105 0.66 2.105 1.395 2.045 1.395 2.045 0.66 1.74 0.66 1.74 0.88 1.695 0.88 1.695 1.395 1.635 1.395 1.635 0.83 1.655 0.83 1.655 0.415 1.61 0.415 1.61 0.295 1.67 0.295 1.67 0.355 1.715 0.355 1.715 0.6 2.02 0.6 2.02 0.235 2.08 0.235 2.08 0.6 2.41 0.6 2.41 0.485 2.43 0.485 2.43 0.235 2.49 0.235 2.49 0.545 2.47 0.545 2.47 0.925 2.515 0.925 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.675 1.34 1.175 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 0.995 0.46 0.995 0.46 0.79 0.58 0.79 0.58 0.615 0.66 0.615 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.039375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.7714285 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.84 1.175 0.28 1.175 0.28 1.11 0.26 1.11 0.26 0.915 0.36 0.915 0.36 1.095 0.76 1.095 0.76 0.915 0.84 0.915 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 1.77 0 1.77 0 1.65 0.375 1.65 0.375 1.275 0.435 1.275 0.435 1.65 1.43 1.65 1.43 1.275 1.49 1.275 1.49 1.65 1.84 1.65 1.84 0.925 1.9 0.925 1.9 1.65 2.25 1.65 2.25 0.925 2.31 0.925 2.31 1.65 2.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 0.06 2.285 0.06 2.285 0.5 2.225 0.5 2.225 0.06 1.875 0.06 1.875 0.5 1.815 0.5 1.815 0.06 1.395 0.06 1.395 0.355 1.335 0.355 1.335 0.06 0.585 0.06 0.585 0.355 0.525 0.355 0.525 0.06 0 0.06 0 -0.06 2.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.555 0.73 1.495 0.73 1.495 0.575 1.16 0.575 1.16 1.18 1 1.18 1 1.24 0.94 1.24 0.94 1.12 1.1 1.12 1.1 0.355 0.835 0.355 0.835 0.235 0.895 0.235 0.895 0.295 1.16 0.295 1.16 0.515 1.555 0.515 ;
      POLYGON 1 1.02 0.94 1.02 0.94 0.815 0.77 0.815 0.77 0.515 0.16 0.515 0.16 1.18 0.18 1.18 0.18 1.3 0.12 1.3 0.12 1.23 0.1 1.23 0.1 0.455 0.225 0.455 0.225 0.32 0.285 0.32 0.285 0.455 0.83 0.455 0.83 0.755 1 0.755 ;
  END
END CLKMX2X6

MACRO CLKMX2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKMX2X8 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.645175 LAYER Metal1 ;
    ANTENNADIFFAREA 2.34975 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.256275 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.41956875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 49.11911025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.325 1.435 3.265 1.435 3.265 1.05 2.915 1.05 2.915 1.435 2.855 1.435 2.855 1.05 2.505 1.05 2.505 1.435 2.445 1.435 2.445 1.05 2.14 1.05 2.14 1.11 2.095 1.11 2.095 1.435 2.035 1.435 2.035 0.99 2.06 0.99 2.06 0.59 2 0.59 2 0.53 2.12 0.53 2.12 0.98 2.14 0.98 2.14 0.99 3.265 0.99 3.265 0.615 2.49 0.615 2.49 0.6 2.415 0.6 2.415 0.54 2.535 0.54 2.535 0.555 2.825 0.555 2.825 0.54 2.945 0.54 2.945 0.555 3.265 0.555 3.265 0.495 3.325 0.495 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 1.19 1.66 1.19 1.66 0.93 1.5 0.93 1.5 0.85 1.74 0.85 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.92556625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.715 0.8 1.085 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.039375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.43809525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.02 0.925 0.96 0.925 0.96 1.245 0.475 1.245 0.475 1.11 0.26 1.11 0.26 0.955 0.535 0.955 0.535 1.185 0.9 1.185 0.9 0.865 1.02 0.865 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 1.77 0 1.77 0 1.65 0.605 1.65 0.605 1.345 0.725 1.345 0.725 1.405 0.665 1.405 0.665 1.65 1.76 1.65 1.76 1.29 1.82 1.29 1.82 1.65 2.24 1.65 2.24 1.15 2.3 1.15 2.3 1.65 2.65 1.65 2.65 1.15 2.71 1.15 2.71 1.65 3.06 1.65 3.06 1.15 3.12 1.15 3.12 1.65 3.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 0.06 3.12 0.06 3.12 0.455 3.06 0.455 3.06 0.06 2.71 0.06 2.71 0.455 2.65 0.455 2.65 0.06 2.295 0.06 2.295 0.455 2.235 0.455 2.235 0.06 1.635 0.06 1.635 0.365 1.695 0.365 1.695 0.425 1.575 0.425 1.575 0.06 0.695 0.06 0.695 0.455 0.635 0.455 0.635 0.06 0 0.06 0 -0.06 3.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.96 0.81 1.9 0.81 1.9 0.75 1.4 0.75 1.4 1.19 1.145 1.19 1.145 1.435 1.085 1.435 1.085 1.13 1.34 1.13 1.34 0.455 1.19 0.455 1.19 0.335 1.25 0.335 1.25 0.395 1.4 0.395 1.4 0.69 1.96 0.69 ;
      POLYGON 1.24 0.695 1.18 0.695 1.18 0.97 1.24 0.97 1.24 1.03 1.12 1.03 1.12 0.615 0.16 0.615 0.16 1.21 0.375 1.21 0.375 1.33 0.315 1.33 0.315 1.27 0.1 1.27 0.1 0.555 0.4 0.555 0.4 0.42 0.46 0.42 0.46 0.555 1.18 0.555 1.18 0.635 1.24 0.635 ;
  END
END CLKMX2X8

MACRO CLKXOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKXOR2X1 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.841925 LAYER Metal1 ;
    ANTENNADIFFAREA 0.8979 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06165 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.65652875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 112.77372275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.14 0.54 0.13 0.54 0.13 1.29 0.07 1.29 0.07 0.54 0.06 0.54 0.06 0.41 0.07 0.41 0.07 0.275 0.13 0.275 0.13 0.41 0.14 0.41 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.58333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.335 0.905 1.275 0.905 1.275 0.875 1.165 0.875 1.165 0.92 1.035 0.92 1.035 0.875 0.9 0.875 0.9 0.97 0.72 0.97 0.72 1.045 0.66 1.045 0.66 0.91 0.84 0.91 0.84 0.815 1.035 0.815 1.035 0.79 1.165 0.79 1.165 0.815 1.275 0.815 1.275 0.785 1.335 0.785 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.9814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.59 0.73 0.45 0.73 0.45 0.885 0.39 0.885 0.39 0.6 0.59 0.6 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.49 0.395 1.49 0.395 1.65 1.125 1.65 1.125 1.17 1.185 1.17 1.185 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.205 0.06 1.205 0.445 1.145 0.445 1.145 0.06 0.335 0.06 0.335 0.395 0.275 0.395 0.275 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.455 1.07 1.39 1.07 1.39 1.195 1.305 1.195 1.305 1.07 1.025 1.07 1.025 1.42 0.85 1.42 0.85 1.36 0.965 1.36 0.965 1.01 1.395 1.01 1.395 0.47 1.35 0.47 1.35 0.35 1.41 0.35 1.41 0.41 1.455 0.41 ;
      POLYGON 1.205 0.715 0.73 0.715 0.73 0.85 0.58 0.85 0.58 1.195 0.52 1.195 0.52 0.79 0.67 0.79 0.67 0.47 0.52 0.47 0.52 0.35 0.58 0.35 0.58 0.41 0.73 0.41 0.73 0.655 1.205 0.655 ;
      POLYGON 0.895 0.445 0.835 0.445 0.835 0.265 0.455 0.265 0.455 0.54 0.29 0.54 0.29 1.33 0.69 1.33 0.69 1.2 0.725 1.2 0.725 1.14 0.785 1.14 0.785 1.26 0.75 1.26 0.75 1.39 0.23 1.39 0.23 0.48 0.395 0.48 0.395 0.205 0.895 0.205 ;
  END
END CLKXOR2X1

MACRO CLKXOR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKXOR2X2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0182 LAYER Metal1 ;
    ANTENNADIFFAREA 1.164775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0909 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.20132025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 91.320132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.435 0.555 0.34 0.555 0.34 1.155 0.435 1.155 0.435 1.275 0.375 1.275 0.375 1.215 0.28 1.215 0.28 0.73 0.26 0.73 0.26 0.6 0.28 0.6 0.28 0.495 0.375 0.495 0.375 0.435 0.435 0.435 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.45370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.785 0.875 1.565 0.875 1.565 0.895 1.435 0.895 1.435 0.885 1.06 0.885 1.06 0.825 1.335 0.825 1.335 0.815 1.785 0.815 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.195 0.72 1.195 0.72 0.895 0.6 0.895 0.6 0.815 0.8 0.815 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.12 1.65 0.12 0.985 0.18 0.985 0.18 1.65 0.58 1.65 0.58 1.54 0.7 1.54 0.7 1.65 1.52 1.65 1.52 1.17 1.58 1.17 1.58 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.625 0.06 1.625 0.55 1.565 0.55 1.565 0.06 0.64 0.06 0.64 0.52 0.58 0.52 0.58 0.06 0.18 0.06 0.18 0.52 0.12 0.52 0.12 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.945 1.07 1.785 1.07 1.785 1.195 1.725 1.195 1.725 1.07 1.42 1.07 1.42 1.42 1.22 1.42 1.22 1.36 1.36 1.36 1.36 1.01 1.885 1.01 1.885 0.575 1.77 0.575 1.77 0.455 1.83 0.455 1.83 0.515 1.945 0.515 ;
      POLYGON 1.625 0.715 0.96 0.715 0.96 1.195 0.9 1.195 0.9 0.485 1.02 0.485 1.02 0.545 0.96 0.545 0.96 0.655 1.625 0.655 ;
      POLYGON 1.315 0.55 1.255 0.55 1.255 0.385 0.8 0.385 0.8 0.715 0.5 0.715 0.5 0.995 0.62 0.995 0.62 1.295 1.06 1.295 1.06 1.2 1.165 1.2 1.165 1.14 1.225 1.14 1.225 1.26 1.12 1.26 1.12 1.355 0.56 1.355 0.56 1.055 0.44 1.055 0.44 0.655 0.74 0.655 0.74 0.325 1.315 0.325 ;
  END
END CLKXOR2X2

MACRO CLKXOR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKXOR2X4 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.43815 LAYER Metal1 ;
    ANTENNADIFFAREA 1.6488 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.16335 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.8041015 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 70.1928375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.745 0.415 0.7 0.415 0.7 0.575 0.32 0.575 0.32 0.79 0.34 0.79 0.34 0.9 0.7 0.9 0.7 1.155 0.745 1.155 0.745 1.275 0.685 1.275 0.685 1.215 0.64 1.215 0.64 0.96 0.335 0.96 0.335 1.29 0.26 1.29 0.26 0.435 0.335 0.435 0.335 0.515 0.64 0.515 0.64 0.355 0.685 0.355 0.685 0.295 0.745 0.295 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.039375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.6761905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.34 0.92 2.26 0.92 2.26 0.695 1.9 0.695 1.9 0.615 2.34 0.615 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.32 0.755 1.165 0.755 1.165 0.895 0.96 0.895 0.96 0.675 1.32 0.675 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.9 0.13 0.9 0.13 1.65 0.48 1.65 0.48 1.06 0.54 1.06 0.54 1.65 0.89 1.65 0.89 1.275 1.01 1.275 1.01 1.335 0.95 1.335 0.95 1.65 2.175 1.65 2.175 1.155 2.235 1.155 2.235 1.65 2.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 0.06 2.235 0.06 2.235 0.355 2.175 0.355 2.175 0.06 0.95 0.06 0.95 0.415 0.89 0.415 0.89 0.06 0.54 0.06 0.54 0.415 0.48 0.415 0.48 0.06 0.13 0.06 0.13 0.415 0.07 0.415 0.07 0.06 0 0.06 0 -0.06 2.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.5 1.12 2.44 1.12 2.44 1.18 2.38 1.18 2.38 1.06 2.44 1.06 2.44 0.515 1.8 0.515 1.8 0.795 2 0.795 2 0.855 1.74 0.855 1.74 0.63 1.58 0.63 1.58 0.51 1.64 0.51 1.64 0.57 1.74 0.57 1.74 0.455 2.38 0.455 2.38 0.26 2.44 0.26 2.44 0.455 2.5 0.455 ;
      POLYGON 2.16 1.015 1.48 1.015 1.48 1.085 1.42 1.085 1.42 0.35 1.54 0.35 1.54 0.41 1.48 0.41 1.48 0.955 2.1 0.955 2.1 0.795 2.16 0.795 ;
      POLYGON 1.905 1.245 1.11 1.245 1.11 1.175 0.845 1.175 0.845 1.055 0.8 1.055 0.8 0.735 0.59 0.735 0.59 0.675 0.8 0.675 0.8 0.515 1.26 0.515 1.26 0.19 1.87 0.19 1.87 0.355 1.81 0.355 1.81 0.25 1.32 0.25 1.32 0.575 0.86 0.575 0.86 0.995 0.905 0.995 0.905 1.115 1.17 1.115 1.17 1.185 1.845 1.185 1.845 1.125 1.905 1.125 ;
  END
END CLKXOR2X4

MACRO CLKXOR2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN CLKXOR2X8 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.809125 LAYER Metal1 ;
    ANTENNADIFFAREA 2.2778 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.27945 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.47387725 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 50.9178745 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.575 0.54 1.485 0.54 1.485 0.555 0.34 0.555 0.34 0.73 0.32 0.73 0.32 0.915 1.55 0.915 1.55 1.36 1.49 1.36 1.49 0.975 1.14 0.975 1.14 1.36 1.08 1.36 1.08 0.975 0.73 0.975 0.73 1.36 0.67 1.36 0.67 0.975 0.32 0.975 0.32 1.36 0.26 1.36 0.26 0.555 0.255 0.555 0.255 0.435 0.315 0.435 0.315 0.495 0.635 0.495 0.635 0.48 0.755 0.48 0.755 0.495 1.045 0.495 1.045 0.48 1.165 0.48 1.165 0.495 1.44 0.495 1.44 0.48 1.575 0.48 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.039375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.86666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.18 0.87 3.14 0.87 3.14 0.92 3.06 0.92 3.06 0.69 2.72 0.69 2.72 0.61 3.14 0.61 3.14 0.79 3.18 0.79 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.03 1.01 1.95 1.01 1.95 0.745 1.835 0.745 1.835 0.625 2.03 0.625 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 1.77 0 1.77 0 1.65 0.465 1.65 0.465 1.075 0.525 1.075 0.525 1.65 0.875 1.65 0.875 1.075 0.935 1.075 0.935 1.65 1.285 1.65 1.285 1.075 1.345 1.075 1.345 1.65 1.665 1.65 1.665 1.27 1.785 1.27 1.785 1.33 1.725 1.33 1.725 1.65 2.92 1.65 2.92 1.14 2.98 1.14 2.98 1.65 3.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 0.06 3.055 0.06 3.055 0.35 2.995 0.35 2.995 0.06 1.72 0.06 1.72 0.305 1.78 0.305 1.78 0.365 1.66 0.365 1.66 0.06 1.34 0.06 1.34 0.395 1.28 0.395 1.28 0.06 0.93 0.06 0.93 0.395 0.87 0.395 0.87 0.06 0.52 0.06 0.52 0.395 0.46 0.395 0.46 0.06 0 0.06 0 -0.06 3.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.34 1.08 3.215 1.08 3.215 1.14 3.155 1.14 3.155 1.02 3.28 1.02 3.28 0.51 2.61 0.51 2.61 0.79 2.67 0.79 2.67 0.85 2.55 0.85 2.55 0.665 2.375 0.665 2.375 0.725 2.315 0.725 2.315 0.605 2.55 0.605 2.55 0.45 3.27 0.45 3.27 0.255 3.34 0.255 ;
      POLYGON 2.915 1.01 2.215 1.01 2.215 1.07 2.155 1.07 2.155 0.345 2.275 0.345 2.275 0.405 2.215 0.405 2.215 0.95 2.855 0.95 2.855 0.79 2.915 0.79 ;
      POLYGON 2.61 1.23 1.885 1.23 1.885 1.17 1.675 1.17 1.675 0.715 1.125 0.715 1.125 0.655 1.675 0.655 1.675 0.465 1.88 0.465 1.88 0.185 2.505 0.185 2.505 0.35 2.445 0.35 2.445 0.245 1.94 0.245 1.94 0.525 1.735 0.525 1.735 1.11 1.945 1.11 1.945 1.17 2.55 1.17 2.55 1.11 2.61 1.11 ;
  END
END CLKXOR2X8

MACRO DECAP2
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN DECAP2 0 0 ;
  SIZE 0.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.4 1.77 0 1.77 0 1.65 0.08 1.65 0.08 0.735 0.05 0.735 0.05 0.675 0.17 0.675 0.17 0.735 0.14 0.735 0.14 1.08 0.27 1.08 0.27 0.95 0.33 0.95 0.33 1.36 0.27 1.36 0.27 1.14 0.14 1.14 0.14 1.65 0.4 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.4 0.06 0.33 0.06 0.33 0.875 0.27 0.875 0.27 0.51 0.13 0.51 0.13 0.6 0.07 0.6 0.07 0.35 0.13 0.35 0.13 0.45 0.27 0.45 0.27 0.06 0 0.06 0 -0.06 0.4 -0.06 ;
    END
  END VSS
END DECAP2

MACRO DECAP3
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN DECAP3 0 0 ;
  SIZE 0.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.74 0.04 0.74 0.04 0.68 0.16 0.68 0.16 0.74 0.13 0.74 0.13 1.65 0.47 1.65 0.47 0.95 0.53 0.95 0.53 1.65 0.6 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 0.06 0.53 0.06 0.53 0.82 0.56 0.82 0.56 0.88 0.44 0.88 0.44 0.82 0.47 0.82 0.47 0.06 0.13 0.06 0.13 0.61 0.07 0.61 0.07 0.06 0 0.06 0 -0.06 0.6 -0.06 ;
    END
  END VSS
END DECAP3

MACRO DECAP4
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN DECAP4 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.74 0.04 0.74 0.04 0.68 0.16 0.68 0.16 0.74 0.13 0.74 0.13 1.65 0.67 1.65 0.67 0.95 0.73 0.95 0.73 1.65 0.8 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 0.06 0.73 0.06 0.73 0.82 0.76 0.82 0.76 0.88 0.64 0.88 0.64 0.82 0.67 0.82 0.67 0.06 0.13 0.06 0.13 0.61 0.07 0.61 0.07 0.06 0 0.06 0 -0.06 0.8 -0.06 ;
    END
  END VSS
END DECAP4

MACRO DECAP5
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DECAP5 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.74 0.04 0.74 0.04 0.68 0.16 0.68 0.16 0.74 0.13 0.74 0.13 1.65 0.87 1.65 0.87 0.95 0.93 0.95 0.93 1.65 1 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.93 0.06 0.93 0.82 0.96 0.82 0.96 0.88 0.84 0.88 0.84 0.82 0.87 0.82 0.87 0.06 0.13 0.06 0.13 0.61 0.07 0.61 0.07 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
  END VSS
END DECAP5

MACRO DECAP6
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN DECAP6 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.74 0.04 0.74 0.04 0.68 0.525 0.68 0.525 0.74 0.13 0.74 0.13 1.65 1.07 1.65 1.07 0.95 1.13 0.95 1.13 1.65 1.2 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 1.13 0.06 1.13 0.82 1.16 0.82 1.16 0.88 0.68 0.88 0.68 0.82 1.07 0.82 1.07 0.06 0.13 0.06 0.13 0.61 0.07 0.61 0.07 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
  END VSS
END DECAP6

MACRO DECAP7
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN DECAP7 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.74 0.04 0.74 0.04 0.68 0.64 0.68 0.64 0.74 0.13 0.74 0.13 1.65 1.27 1.65 1.27 0.95 1.33 0.95 1.33 1.65 1.4 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 1.33 0.06 1.33 0.82 1.36 0.82 1.36 0.88 0.76 0.88 0.76 0.82 1.27 0.82 1.27 0.06 0.13 0.06 0.13 0.61 0.07 0.61 0.07 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
  END VSS
END DECAP7

MACRO DECAP8
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN DECAP8 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.74 0.04 0.74 0.04 0.68 0.77 0.68 0.77 0.74 0.13 0.74 0.13 1.65 1.47 1.65 1.47 0.95 1.53 0.95 1.53 1.65 1.6 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.53 0.06 1.53 0.82 1.56 0.82 1.56 0.88 0.83 0.88 0.83 0.82 1.47 0.82 1.47 0.06 0.13 0.06 0.13 0.61 0.07 0.61 0.07 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
  END VSS
END DECAP8

MACRO DECAP9
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN DECAP9 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.74 0.04 0.74 0.04 0.68 0.885 0.68 0.885 0.74 0.13 0.74 0.13 1.65 1.67 1.65 1.67 0.95 1.73 0.95 1.73 1.65 1.8 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.73 0.06 1.73 0.82 1.76 0.82 1.76 0.88 0.93 0.88 0.93 0.82 1.67 0.82 1.67 0.06 0.13 0.06 0.13 0.61 0.07 0.61 0.07 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
  END VSS
END DECAP9

MACRO DECAP10
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN DECAP10 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.74 0.04 0.74 0.04 0.68 0.885 0.68 0.885 0.74 0.13 0.74 0.13 1.65 1.87 1.65 1.87 0.95 1.93 0.95 1.93 1.65 2 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.93 0.06 1.93 0.82 1.96 0.82 1.96 0.88 1 0.88 1 0.82 1.87 0.82 1.87 0.06 0.13 0.06 0.13 0.61 0.07 0.61 0.07 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
  END VSS
END DECAP10

MACRO DFF2RX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFF2RX1 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.045 0.77 4.225 0.92 ;
    END
  END CK
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5614 LAYER Metal1 ;
    ANTENNADIFFAREA 6.234075 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4248 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.737759 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.03531075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.75 1.18 0.69 1.18 0.69 0.765 0.65 0.765 0.65 0.4 0.75 0.4 ;
    END
  END Q1
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5614 LAYER Metal1 ;
    ANTENNADIFFAREA 6.266525 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4248 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.737759 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.03531075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.05 0.4 0.14 1.155 ;
    END
  END Q1N
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.395 0.625 3.54 0.905 ;
    END
  END D1
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0648 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 26.3425925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.78 1.48 1.22 1.48 1.22 1.42 3.06 1.42 3.06 1.385 3.345 1.385 3.345 1.42 4.655 1.42 4.655 1.385 4.94 1.385 4.94 1.42 6.78 1.42 ;
    END
  END RN
  PIN Q2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5614 LAYER Metal1 ;
    ANTENNADIFFAREA 5.884175 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4248 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.737759 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.03531075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.35 0.765 7.31 0.765 7.31 1.18 7.25 1.18 7.25 0.4 7.35 0.4 ;
    END
  END Q2
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5614 LAYER Metal1 ;
    ANTENNADIFFAREA 6.86445 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4248 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.737759 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.03531075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.86 0.4 7.95 1.155 ;
    END
  END Q2N
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.46 0.625 4.605 0.905 ;
    END
  END D2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.54 0.395 1.54 0.395 1.65 0.855 1.65 0.855 1.54 0.975 1.54 0.975 1.65 1.42 1.65 1.42 1.54 1.54 1.54 1.54 1.65 2.125 1.65 2.125 1.54 2.245 1.54 2.245 1.65 2.52 1.65 2.52 1.54 2.645 1.54 2.645 1.65 3.435 1.65 3.435 1.54 3.555 1.54 3.555 1.65 3.93 1.65 3.93 1.54 4.05 1.54 4.05 1.65 4.445 1.65 4.445 1.54 4.565 1.54 4.565 1.65 5.355 1.65 5.355 1.54 5.48 1.54 5.48 1.65 5.755 1.65 5.755 1.54 5.875 1.54 5.875 1.65 6.46 1.65 6.46 1.54 6.58 1.54 6.58 1.65 7.025 1.65 7.025 1.54 7.145 1.54 7.145 1.65 7.605 1.65 7.605 1.54 7.725 1.54 7.725 1.65 8 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 0.06 7.7 0.06 7.7 0.17 7.58 0.17 7.58 0.06 7.175 0.06 7.175 0.17 7.055 0.17 7.055 0.06 6.655 0.06 6.655 0.17 6.52 0.17 6.52 0.06 5.8 0.06 5.8 0.17 5.68 0.17 5.68 0.06 4.57 0.06 4.57 0.17 4.45 0.17 4.45 0.165 4.445 0.165 4.445 0.06 4.05 0.06 4.05 0.17 3.925 0.17 3.925 0.06 3.555 0.06 3.555 0.165 3.55 0.165 3.55 0.17 3.43 0.17 3.43 0.06 2.32 0.06 2.32 0.17 2.2 0.17 2.2 0.06 1.48 0.06 1.48 0.17 1.345 0.17 1.345 0.06 0.945 0.06 0.945 0.17 0.825 0.17 0.825 0.06 0.42 0.06 0.42 0.17 0.3 0.17 0.3 0.06 0 0.06 0 -0.06 8 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.78 0.86 7.72 0.86 7.72 0.83 7.53 0.83 7.53 1.02 7.47 1.02 7.47 0.54 7.53 0.54 7.53 0.77 7.72 0.77 7.72 0.74 7.78 0.74 ;
      POLYGON 7.185 0.83 7 0.83 7 1.12 6.49 1.12 6.49 0.765 6.55 0.765 6.55 1.06 6.94 1.06 6.94 0.49 6.795 0.49 6.795 0.43 7 0.43 7 0.77 7.185 0.77 ;
      POLYGON 6.85 0.715 6.79 0.715 6.79 0.685 6.41 0.685 6.41 1.025 6.26 1.025 6.26 1.115 6.2 1.115 6.2 0.965 6.35 0.965 6.35 0.47 6.27 0.47 6.27 0.5 6.21 0.5 6.21 0.375 6.27 0.375 6.27 0.41 6.41 0.41 6.41 0.625 6.79 0.625 6.79 0.595 6.85 0.595 ;
      POLYGON 6.795 0.3 6.13 0.3 6.13 0.615 6.29 0.615 6.29 0.885 6.23 0.885 6.23 0.675 6.07 0.675 6.07 0.3 5.365 0.3 5.365 0.39 5.305 0.39 5.305 0.3 4.855 0.3 4.855 0.855 4.795 0.855 4.795 0.3 4.54 0.3 4.54 0.325 4.445 0.325 4.445 0.3 3.8 0.3 3.8 1.1 3.66 1.1 3.66 0.77 3.74 0.77 3.74 0.3 3.555 0.3 3.555 0.325 3.46 0.325 3.46 0.3 3.205 0.3 3.205 0.855 3.145 0.855 3.145 0.3 2.695 0.3 2.695 0.39 2.635 0.39 2.635 0.3 1.93 0.3 1.93 0.675 1.77 0.675 1.77 0.885 1.71 0.885 1.71 0.615 1.87 0.615 1.87 0.3 1.205 0.3 1.205 0.24 1.87 0.24 1.87 0.185 1.93 0.185 1.93 0.24 6.07 0.24 6.07 0.185 6.13 0.185 6.13 0.24 6.795 0.24 ;
      POLYGON 6.78 1.36 5.03 1.36 5.03 1.3 4.575 1.3 4.575 1.36 3.425 1.36 3.425 1.3 2.97 1.3 2.97 1.36 1.22 1.36 1.22 1.3 2.88 1.3 2.88 1.24 3.425 1.24 3.425 1.195 3.54 1.195 3.54 1.3 3.9 1.3 3.9 0.895 3.86 0.895 3.86 0.495 3.96 0.495 3.96 0.625 4.165 0.625 4.165 0.505 4.225 0.505 4.225 0.705 3.96 0.705 3.96 1.005 4.255 1.005 4.255 1.065 3.96 1.065 3.96 1.3 4.46 1.3 4.46 1.195 4.575 1.195 4.575 1.24 5.12 1.24 5.12 1.3 6.78 1.3 ;
      POLYGON 6.01 1.09 5.95 1.09 5.95 0.71 5.38 0.71 5.38 0.65 5.95 0.65 5.95 0.38 6.01 0.38 ;
      POLYGON 5.87 0.895 5.81 0.895 5.81 0.87 4.975 0.87 4.975 1.15 4.915 1.15 4.915 0.81 5.145 0.81 5.145 0.46 5.205 0.46 5.205 0.81 5.81 0.81 5.81 0.775 5.87 0.775 ;
      RECT 5.085 1.04 5.64 1.1 ;
      RECT 4.665 0.46 4.725 1.14 ;
      RECT 3.275 0.46 3.335 1.14 ;
      POLYGON 3.085 1.15 3.025 1.15 3.025 0.87 2.19 0.87 2.19 0.895 2.13 0.895 2.13 0.775 2.19 0.775 2.19 0.81 2.795 0.81 2.795 0.46 2.855 0.46 2.855 0.81 3.085 0.81 ;
      RECT 2.36 1.04 2.915 1.1 ;
      POLYGON 2.62 0.71 2.05 0.71 2.05 1.09 1.99 1.09 1.99 0.38 2.05 0.38 2.05 0.65 2.62 0.65 ;
      POLYGON 1.8 1.115 1.74 1.115 1.74 1.025 1.59 1.025 1.59 0.685 1.21 0.685 1.21 0.715 1.15 0.715 1.15 0.595 1.21 0.595 1.21 0.625 1.59 0.625 1.59 0.41 1.73 0.41 1.73 0.375 1.79 0.375 1.79 0.5 1.73 0.5 1.73 0.47 1.65 0.47 1.65 0.965 1.8 0.965 ;
      POLYGON 1.51 1.12 1 1.12 1 0.83 0.815 0.83 0.815 0.77 1 0.77 1 0.43 1.205 0.43 1.205 0.49 1.06 0.49 1.06 1.06 1.45 1.06 1.45 0.765 1.51 0.765 ;
      POLYGON 0.53 1.02 0.47 1.02 0.47 0.83 0.28 0.83 0.28 0.86 0.22 0.86 0.22 0.74 0.28 0.74 0.28 0.77 0.47 0.77 0.47 0.54 0.53 0.54 ;
  END
END DFF2RX1

MACRO DFF2RX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFF2RX2 0 0 ;
  SIZE 8.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8656 LAYER Metal1 ;
    ANTENNADIFFAREA 7.37785 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.55575 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.75501575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 63.96221325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.46 0.4 8.55 1.18 ;
    END
  END Q2N
  PIN Q2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8656 LAYER Metal1 ;
    ANTENNADIFFAREA 7.6445 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.55575 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.75501575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 63.96221325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.75 0.755 7.71 0.755 7.71 1.18 7.65 1.18 7.65 0.4 7.75 0.4 ;
    END
  END Q2
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.86 0.625 5.005 0.905 ;
    END
  END D2
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.07875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 21.6761905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.18 1.48 1.62 1.48 1.62 1.42 3.46 1.42 3.46 1.385 3.745 1.385 3.745 1.42 5.055 1.42 5.055 1.385 5.34 1.385 5.34 1.42 7.18 1.42 ;
    END
  END RN
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8656 LAYER Metal1 ;
    ANTENNADIFFAREA 7.39765 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.55575 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.75501575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 63.96221325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 0.4 0.34 1.18 ;
    END
  END Q1N
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8656 LAYER Metal1 ;
    ANTENNADIFFAREA 7.355425 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.55575 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.75501575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 63.96221325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.15 1.18 1.09 1.18 1.09 0.755 1.05 0.755 1.05 0.4 1.15 0.4 ;
    END
  END Q1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.795 0.625 3.94 0.905 ;
    END
  END D1
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.445 0.77 4.625 0.92 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.8 1.77 0 1.77 0 1.65 0.055 1.65 0.055 1.54 0.175 1.54 0.175 1.65 0.475 1.65 0.475 1.54 0.595 1.54 0.595 1.65 0.82 1.65 0.82 1.54 0.94 1.54 0.94 1.65 1.255 1.65 1.255 1.54 1.375 1.54 1.375 1.65 1.82 1.65 1.82 1.54 1.94 1.54 1.94 1.65 2.525 1.65 2.525 1.54 2.645 1.54 2.645 1.65 2.92 1.65 2.92 1.54 3.045 1.54 3.045 1.65 3.835 1.65 3.835 1.54 3.955 1.54 3.955 1.65 4.33 1.65 4.33 1.54 4.45 1.54 4.45 1.65 4.845 1.65 4.845 1.54 4.965 1.54 4.965 1.65 5.755 1.65 5.755 1.54 5.88 1.54 5.88 1.65 6.155 1.65 6.155 1.54 6.275 1.54 6.275 1.65 6.86 1.65 6.86 1.54 6.98 1.54 6.98 1.65 7.425 1.65 7.425 1.54 7.545 1.54 7.545 1.65 7.86 1.65 7.86 1.54 7.98 1.54 7.98 1.65 8.205 1.65 8.205 1.54 8.325 1.54 8.325 1.65 8.625 1.65 8.625 1.54 8.745 1.54 8.745 1.65 8.8 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.8 0.06 8.745 0.06 8.745 0.17 8.625 0.17 8.625 0.06 8.3 0.06 8.3 0.17 8.18 0.17 8.18 0.06 7.945 0.06 7.945 0.17 7.825 0.17 7.825 0.06 7.575 0.06 7.575 0.17 7.455 0.17 7.455 0.06 7.055 0.06 7.055 0.17 6.935 0.17 6.935 0.165 6.92 0.165 6.92 0.06 6.2 0.06 6.2 0.17 6.08 0.17 6.08 0.06 4.97 0.06 4.97 0.17 4.845 0.17 4.845 0.06 4.45 0.06 4.45 0.17 4.325 0.17 4.325 0.06 3.955 0.06 3.955 0.17 3.83 0.17 3.83 0.06 2.72 0.06 2.72 0.17 2.6 0.17 2.6 0.06 1.88 0.06 1.88 0.165 1.865 0.165 1.865 0.17 1.745 0.17 1.745 0.06 1.345 0.06 1.345 0.17 1.225 0.17 1.225 0.06 0.975 0.06 0.975 0.17 0.855 0.17 0.855 0.06 0.62 0.06 0.62 0.17 0.5 0.17 0.5 0.06 0.175 0.06 0.175 0.17 0.055 0.17 0.055 0.06 0 0.06 0 -0.06 8.8 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 8.38 0.86 8.32 0.86 8.32 0.83 8.13 0.83 8.13 1.02 8.07 1.02 8.07 0.54 8.13 0.54 8.13 0.77 8.32 0.77 8.32 0.74 8.38 0.74 ;
      POLYGON 7.585 0.83 7.45 0.83 7.45 1.12 6.89 1.12 6.89 0.765 6.95 0.765 6.95 1.06 7.39 1.06 7.39 0.49 7.195 0.49 7.195 0.43 7.45 0.43 7.45 0.77 7.585 0.77 ;
      POLYGON 7.285 0.7 6.81 0.7 6.81 1.025 6.66 1.025 6.66 1.115 6.6 1.115 6.6 0.965 6.75 0.965 6.75 0.47 6.67 0.47 6.67 0.5 6.61 0.5 6.61 0.375 6.67 0.375 6.67 0.41 6.81 0.41 6.81 0.64 7.285 0.64 ;
      POLYGON 7.195 0.3 6.53 0.3 6.53 0.615 6.69 0.615 6.69 0.885 6.63 0.885 6.63 0.675 6.47 0.675 6.47 0.3 5.765 0.3 5.765 0.39 5.705 0.39 5.705 0.3 5.255 0.3 5.255 0.855 5.195 0.855 5.195 0.3 4.94 0.3 4.94 0.325 4.845 0.325 4.845 0.3 4.2 0.3 4.2 1.1 4.06 1.1 4.06 0.77 4.14 0.77 4.14 0.3 3.955 0.3 3.955 0.325 3.86 0.325 3.86 0.3 3.605 0.3 3.605 0.855 3.545 0.855 3.545 0.3 3.095 0.3 3.095 0.39 3.035 0.39 3.035 0.3 2.33 0.3 2.33 0.675 2.17 0.675 2.17 0.885 2.11 0.885 2.11 0.615 2.27 0.615 2.27 0.3 1.605 0.3 1.605 0.24 2.27 0.24 2.27 0.185 2.33 0.185 2.33 0.24 6.47 0.24 6.47 0.185 6.53 0.185 6.53 0.24 7.195 0.24 ;
      POLYGON 7.18 1.36 5.43 1.36 5.43 1.3 4.975 1.3 4.975 1.36 3.825 1.36 3.825 1.3 3.37 1.3 3.37 1.36 1.62 1.36 1.62 1.3 3.28 1.3 3.28 1.24 3.825 1.24 3.825 1.195 3.94 1.195 3.94 1.3 4.3 1.3 4.3 0.895 4.26 0.895 4.26 0.495 4.36 0.495 4.36 0.625 4.565 0.625 4.565 0.505 4.625 0.505 4.625 0.705 4.36 0.705 4.36 1.005 4.655 1.005 4.655 1.065 4.36 1.065 4.36 1.3 4.86 1.3 4.86 1.195 4.975 1.195 4.975 1.24 5.52 1.24 5.52 1.3 7.18 1.3 ;
      POLYGON 6.41 1.09 6.35 1.09 6.35 0.71 5.78 0.71 5.78 0.65 6.35 0.65 6.35 0.38 6.41 0.38 ;
      POLYGON 6.27 0.895 6.21 0.895 6.21 0.87 5.375 0.87 5.375 1.15 5.315 1.15 5.315 0.81 5.545 0.81 5.545 0.46 5.605 0.46 5.605 0.81 6.21 0.81 6.21 0.775 6.27 0.775 ;
      RECT 5.485 1.04 6.04 1.1 ;
      RECT 5.065 0.46 5.125 1.14 ;
      RECT 3.675 0.46 3.735 1.14 ;
      POLYGON 3.485 1.15 3.425 1.15 3.425 0.87 2.59 0.87 2.59 0.895 2.53 0.895 2.53 0.775 2.59 0.775 2.59 0.81 3.195 0.81 3.195 0.46 3.255 0.46 3.255 0.81 3.485 0.81 ;
      RECT 2.76 1.04 3.315 1.1 ;
      POLYGON 3.02 0.71 2.45 0.71 2.45 1.09 2.39 1.09 2.39 0.38 2.45 0.38 2.45 0.65 3.02 0.65 ;
      POLYGON 2.2 1.115 2.14 1.115 2.14 1.025 1.99 1.025 1.99 0.7 1.515 0.7 1.515 0.64 1.99 0.64 1.99 0.41 2.13 0.41 2.13 0.375 2.19 0.375 2.19 0.5 2.13 0.5 2.13 0.47 2.05 0.47 2.05 0.965 2.2 0.965 ;
      POLYGON 1.91 1.12 1.35 1.12 1.35 0.83 1.215 0.83 1.215 0.77 1.35 0.77 1.35 0.43 1.605 0.43 1.605 0.49 1.41 0.49 1.41 1.06 1.85 1.06 1.85 0.765 1.91 0.765 ;
      POLYGON 0.73 1.02 0.67 1.02 0.67 0.83 0.48 0.83 0.48 0.86 0.42 0.86 0.42 0.74 0.48 0.74 0.48 0.77 0.67 0.77 0.67 0.54 0.73 0.54 ;
  END
END DFF2RX2

MACRO DFF2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFF2X1 0 0 ;
  SIZE 7.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.645 0.77 3.825 0.92 ;
    END
  END CK
  PIN Q2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1411 LAYER Metal1 ;
    ANTENNADIFFAREA 5.67385 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4248 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.74835225 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 71.0805085 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.545 1.29 6.41 1.29 6.41 0.41 6.47 0.41 6.47 0.9 6.545 0.9 ;
    END
  END Q2
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.25925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.06 0.77 4.185 1.145 ;
    END
  END D2
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1411 LAYER Metal1 ;
    ANTENNADIFFAREA 5.67385 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4248 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.74835225 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 71.0805085 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.14 0.93 7.11 0.93 7.11 1.29 7.05 1.29 7.05 0.41 7.11 0.41 7.11 0.6 7.14 0.6 ;
    END
  END Q2N
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1411 LAYER Metal1 ;
    ANTENNADIFFAREA 5.67385 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4248 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.74835225 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 71.0805085 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.79 1.29 0.655 1.29 0.655 0.9 0.73 0.9 0.73 0.41 0.79 0.41 ;
    END
  END Q1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.25925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.015 0.77 3.14 1.145 ;
    END
  END D1
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.1411 LAYER Metal1 ;
    ANTENNADIFFAREA 5.67385 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4248 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.74835225 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 71.0805085 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.29 0.09 1.29 0.09 0.93 0.06 0.93 0.06 0.6 0.09 0.6 0.09 0.41 0.15 0.41 ;
    END
  END Q1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 1.77 0 1.77 0 1.65 0.245 1.65 0.245 1.54 0.365 1.54 0.365 1.65 0.935 1.65 0.935 1.54 1.055 1.54 1.055 1.65 1.28 1.65 1.28 1.54 1.4 1.54 1.4 1.65 2.1 1.65 2.1 1.54 2.22 1.54 2.22 1.65 3.015 1.65 3.015 1.54 3.135 1.54 3.135 1.65 3.53 1.65 3.53 1.54 3.65 1.54 3.65 1.65 4.065 1.65 4.065 1.54 4.185 1.54 4.185 1.65 4.98 1.65 4.98 1.54 5.1 1.54 5.1 1.65 5.8 1.65 5.8 1.54 5.92 1.54 5.92 1.65 6.145 1.65 6.145 1.54 6.265 1.54 6.265 1.65 6.835 1.65 6.835 1.54 6.955 1.54 6.955 1.65 7.2 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 0.06 6.955 0.06 6.955 0.17 6.835 0.17 6.835 0.06 6.265 0.06 6.265 0.17 6.145 0.17 6.145 0.06 5.895 0.06 5.895 0.17 5.775 0.17 5.775 0.06 4.985 0.06 4.985 0.17 4.865 0.17 4.865 0.06 4.185 0.06 4.185 0.17 4.065 0.17 4.065 0.06 3.65 0.06 3.65 0.17 3.525 0.17 3.525 0.06 3.135 0.06 3.135 0.17 3.015 0.17 3.015 0.06 2.335 0.06 2.335 0.17 2.215 0.17 2.215 0.06 1.425 0.06 1.425 0.17 1.305 0.17 1.305 0.06 1.055 0.06 1.055 0.17 0.935 0.17 0.935 0.06 0.365 0.06 0.365 0.17 0.245 0.17 0.245 0.06 0 0.06 0 -0.06 7.2 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.97 0.82 6.91 0.82 6.91 0.79 6.69 0.79 6.69 1.02 6.63 1.02 6.63 0.54 6.69 0.54 6.69 0.7 6.97 0.7 ;
      POLYGON 6.31 0.82 6.25 0.82 6.25 0.68 6.07 0.68 6.07 1.21 6.01 1.21 6.01 0.765 5.825 0.765 5.825 0.825 5.765 0.825 5.765 0.705 6.01 0.705 6.01 0.47 6.07 0.47 6.07 0.62 6.31 0.62 ;
      POLYGON 5.945 0.985 5.705 0.985 5.705 1.18 5.435 1.18 5.435 1.12 5.645 1.12 5.645 0.6 5.445 0.6 5.445 0.54 5.705 0.54 5.705 0.925 5.885 0.925 5.885 0.865 5.945 0.865 ;
      POLYGON 5.69 0.31 5.375 0.31 5.375 0.79 5.545 0.79 5.545 1.035 5.485 1.035 5.485 0.85 5.315 0.85 5.315 0.31 4.68 0.31 4.68 0.44 4.62 0.44 4.62 0.345 4.38 0.345 4.38 0.31 3.4 0.31 3.4 1.1 3.26 1.1 3.26 0.77 3.34 0.77 3.34 0.31 2.82 0.31 2.82 0.345 2.58 0.345 2.58 0.44 2.52 0.44 2.52 0.31 1.885 0.31 1.885 0.85 1.715 0.85 1.715 1.035 1.655 1.035 1.655 0.79 1.825 0.79 1.825 0.31 1.51 0.31 1.51 0.25 2.52 0.25 2.52 0.22 2.82 0.22 2.82 0.25 4.38 0.25 4.38 0.22 4.68 0.22 4.68 0.25 5.69 0.25 ;
      POLYGON 5.545 1.48 1.655 1.48 1.655 1.42 1.825 1.42 1.825 0.93 1.885 0.93 1.885 1.42 2.665 1.42 2.665 0.695 2.725 0.695 2.725 1.385 3 1.385 3 1.42 3.46 1.42 3.46 0.495 3.56 0.495 3.56 0.625 3.765 0.625 3.765 0.505 3.825 0.505 3.825 0.705 3.56 0.705 3.56 1.005 3.855 1.005 3.855 1.065 3.54 1.065 3.54 1.42 4.2 1.42 4.2 1.385 4.475 1.385 4.475 0.695 4.535 0.695 4.535 1.42 5.315 1.42 5.315 0.93 5.375 0.93 5.375 1.42 5.545 1.42 ;
      POLYGON 5.255 1.22 5.195 1.22 5.195 0.785 4.905 0.785 4.905 0.725 5.19 0.725 5.19 0.475 5.255 0.475 ;
      POLYGON 5.08 1.005 5.02 1.005 5.02 0.945 4.835 0.945 4.835 1.18 4.635 1.18 4.635 1.12 4.775 1.12 4.775 0.63 4.555 0.63 4.555 0.51 4.615 0.51 4.615 0.57 4.835 0.57 4.835 0.885 5.08 0.885 ;
      RECT 4.33 0.48 4.39 1.22 ;
      RECT 2.81 0.48 2.87 1.22 ;
      POLYGON 2.645 0.63 2.425 0.63 2.425 1.12 2.565 1.12 2.565 1.18 2.365 1.18 2.365 0.945 2.18 0.945 2.18 1.005 2.12 1.005 2.12 0.885 2.365 0.885 2.365 0.57 2.585 0.57 2.585 0.51 2.645 0.51 ;
      POLYGON 2.295 0.785 2.005 0.785 2.005 1.22 1.945 1.22 1.945 0.475 2.01 0.475 2.01 0.725 2.295 0.725 ;
      POLYGON 1.765 1.18 1.495 1.18 1.495 0.985 1.255 0.985 1.255 0.865 1.315 0.865 1.315 0.925 1.495 0.925 1.495 0.54 1.755 0.54 1.755 0.6 1.555 0.6 1.555 1.12 1.765 1.12 ;
      POLYGON 1.435 0.825 1.375 0.825 1.375 0.765 1.19 0.765 1.19 1.21 1.13 1.21 1.13 0.68 0.95 0.68 0.95 0.82 0.89 0.82 0.89 0.62 1.13 0.62 1.13 0.47 1.19 0.47 1.19 0.705 1.435 0.705 ;
      POLYGON 0.57 1.02 0.51 1.02 0.51 0.79 0.29 0.79 0.29 0.82 0.23 0.82 0.23 0.7 0.51 0.7 0.51 0.54 0.57 0.54 ;
  END
END DFF2X1

MACRO DFF2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFF2X2 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.045 0.77 4.225 0.92 ;
    END
  END CK
  PIN Q2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5302 LAYER Metal1 ;
    ANTENNADIFFAREA 6.726775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.55575 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.151507 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 58.40755725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.02 1.085 6.86 1.085 6.86 1.29 6.8 1.29 6.8 0.9 6.96 0.9 6.96 0.66 6.8 0.66 6.8 0.41 6.86 0.41 6.86 0.595 7.02 0.595 ;
    END
  END Q2
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.25925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.46 0.77 4.585 1.145 ;
    END
  END D2
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5302 LAYER Metal1 ;
    ANTENNADIFFAREA 6.726775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.55575 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.151507 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 58.40755725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.74 0.93 7.67 0.93 7.67 1.29 7.61 1.29 7.61 0.41 7.67 0.41 7.67 0.6 7.74 0.6 ;
    END
  END Q2N
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5302 LAYER Metal1 ;
    ANTENNADIFFAREA 6.726775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.55575 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.151507 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 58.40755725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.66 1.04 0.66 1.04 0.9 1.2 0.9 1.2 1.29 1.14 1.29 1.14 1.085 0.98 1.085 0.98 0.595 1.14 0.595 1.14 0.41 1.2 0.41 ;
    END
  END Q1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.25925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.415 0.77 3.54 1.145 ;
    END
  END D1
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5302 LAYER Metal1 ;
    ANTENNADIFFAREA 6.726775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.55575 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.151507 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 58.40755725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.39 1.29 0.33 1.29 0.33 0.93 0.26 0.93 0.26 0.705 0.255 0.705 0.255 0.625 0.26 0.625 0.26 0.6 0.33 0.6 0.33 0.41 0.39 0.41 ;
    END
  END Q1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 1.77 0 1.77 0 1.65 0.115 1.65 0.115 1.54 0.235 1.54 0.235 1.65 0.485 1.65 0.485 1.54 0.605 1.54 0.605 1.65 0.94 1.65 0.94 1.54 1.06 1.54 1.06 1.65 1.28 1.65 1.28 1.54 1.4 1.54 1.4 1.65 1.735 1.65 1.735 1.54 1.855 1.54 1.855 1.65 2.5 1.65 2.5 1.54 2.62 1.54 2.62 1.65 3.415 1.65 3.415 1.54 3.535 1.54 3.535 1.65 3.93 1.65 3.93 1.54 4.05 1.54 4.05 1.65 4.465 1.65 4.465 1.54 4.585 1.54 4.585 1.65 5.38 1.65 5.38 1.54 5.5 1.54 5.5 1.65 6.145 1.65 6.145 1.54 6.265 1.54 6.265 1.65 6.6 1.65 6.6 1.54 6.72 1.54 6.72 1.65 6.94 1.65 6.94 1.54 7.06 1.54 7.06 1.65 7.395 1.65 7.395 1.54 7.515 1.54 7.515 1.65 7.765 1.65 7.765 1.54 7.885 1.54 7.885 1.65 8 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 0.06 7.885 0.06 7.885 0.17 7.765 0.17 7.765 0.06 7.515 0.06 7.515 0.17 7.395 0.17 7.395 0.06 7.06 0.06 7.06 0.17 6.94 0.17 6.94 0.06 6.72 0.06 6.72 0.17 6.6 0.17 6.6 0.06 6.295 0.06 6.295 0.17 6.175 0.17 6.175 0.06 5.385 0.06 5.385 0.17 5.265 0.17 5.265 0.06 4.585 0.06 4.585 0.17 4.465 0.17 4.465 0.06 4.05 0.06 4.05 0.17 3.925 0.17 3.925 0.06 3.535 0.06 3.535 0.17 3.415 0.17 3.415 0.06 2.735 0.06 2.735 0.17 2.615 0.17 2.615 0.06 1.825 0.06 1.825 0.17 1.705 0.17 1.705 0.06 1.4 0.06 1.4 0.17 1.28 0.17 1.28 0.06 1.06 0.06 1.06 0.17 0.94 0.17 0.94 0.06 0.605 0.06 0.605 0.17 0.485 0.17 0.485 0.06 0.235 0.06 0.235 0.17 0.115 0.17 0.115 0.06 0 0.06 0 -0.06 8 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.53 0.82 7.47 0.82 7.47 0.79 7.25 0.79 7.25 1.02 7.19 1.02 7.19 0.54 7.25 0.54 7.25 0.7 7.53 0.7 ;
      POLYGON 6.895 0.8 6.47 0.8 6.47 1.33 6.41 1.33 6.41 0.765 6.225 0.765 6.225 0.825 6.165 0.825 6.165 0.705 6.41 0.705 6.41 0.41 6.47 0.41 6.47 0.74 6.895 0.74 ;
      POLYGON 6.345 0.985 6.105 0.985 6.105 1.18 5.835 1.18 5.835 1.12 6.045 1.12 6.045 0.6 5.845 0.6 5.845 0.54 6.105 0.54 6.105 0.925 6.285 0.925 6.285 0.865 6.345 0.865 ;
      POLYGON 6.09 0.31 5.775 0.31 5.775 0.79 5.945 0.79 5.945 1.035 5.885 1.035 5.885 0.85 5.715 0.85 5.715 0.31 5.08 0.31 5.08 0.44 5.02 0.44 5.02 0.345 4.78 0.345 4.78 0.31 3.8 0.31 3.8 1.1 3.66 1.1 3.66 0.77 3.74 0.77 3.74 0.31 3.22 0.31 3.22 0.345 2.98 0.345 2.98 0.44 2.92 0.44 2.92 0.31 2.285 0.31 2.285 0.85 2.115 0.85 2.115 1.035 2.055 1.035 2.055 0.79 2.225 0.79 2.225 0.31 1.91 0.31 1.91 0.25 2.92 0.25 2.92 0.22 3.22 0.22 3.22 0.25 4.78 0.25 4.78 0.22 5.08 0.22 5.08 0.25 6.09 0.25 ;
      POLYGON 6.08 1.48 1.92 1.48 1.92 1.42 2.225 1.42 2.225 0.93 2.285 0.93 2.285 1.42 3.065 1.42 3.065 0.695 3.125 0.695 3.125 1.385 3.4 1.385 3.4 1.42 3.86 1.42 3.86 0.495 3.96 0.495 3.96 0.625 4.165 0.625 4.165 0.505 4.225 0.505 4.225 0.705 3.96 0.705 3.96 1.005 4.255 1.005 4.255 1.065 3.94 1.065 3.94 1.42 4.6 1.42 4.6 1.385 4.875 1.385 4.875 0.695 4.935 0.695 4.935 1.42 5.715 1.42 5.715 0.93 5.775 0.93 5.775 1.42 6.08 1.42 ;
      POLYGON 5.655 1.22 5.595 1.22 5.595 0.785 5.305 0.785 5.305 0.725 5.59 0.725 5.59 0.475 5.655 0.475 ;
      POLYGON 5.48 1.005 5.42 1.005 5.42 0.945 5.235 0.945 5.235 1.18 5.035 1.18 5.035 1.12 5.175 1.12 5.175 0.63 4.955 0.63 4.955 0.51 5.015 0.51 5.015 0.57 5.235 0.57 5.235 0.885 5.48 0.885 ;
      RECT 4.73 0.48 4.79 1.22 ;
      RECT 3.21 0.48 3.27 1.22 ;
      POLYGON 3.045 0.63 2.825 0.63 2.825 1.12 2.965 1.12 2.965 1.18 2.765 1.18 2.765 0.945 2.58 0.945 2.58 1.005 2.52 1.005 2.52 0.885 2.765 0.885 2.765 0.57 2.985 0.57 2.985 0.51 3.045 0.51 ;
      POLYGON 2.695 0.785 2.405 0.785 2.405 1.22 2.345 1.22 2.345 0.475 2.41 0.475 2.41 0.725 2.695 0.725 ;
      POLYGON 2.165 1.18 1.895 1.18 1.895 0.985 1.655 0.985 1.655 0.865 1.715 0.865 1.715 0.925 1.895 0.925 1.895 0.54 2.155 0.54 2.155 0.6 1.955 0.6 1.955 1.12 2.165 1.12 ;
      POLYGON 1.835 0.825 1.775 0.825 1.775 0.765 1.59 0.765 1.59 1.33 1.53 1.33 1.53 0.8 1.105 0.8 1.105 0.74 1.53 0.74 1.53 0.41 1.59 0.41 1.59 0.705 1.835 0.705 ;
      POLYGON 0.81 1.02 0.75 1.02 0.75 0.79 0.53 0.79 0.53 0.82 0.47 0.82 0.47 0.7 0.75 0.7 0.75 0.54 0.81 0.54 ;
  END
END DFF2X2

MACRO DFF4RX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFF4RX1 0 0 ;
  SIZE 15.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.91405 LAYER Metal1 ;
    ANTENNADIFFAREA 14.03425 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8334 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.69600425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.6299495 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.55 0.765 14.51 0.765 14.51 1.18 14.45 1.18 14.45 0.4 14.55 0.4 ;
    END
  END Q4
  PIN Q4N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.91405 LAYER Metal1 ;
    ANTENNADIFFAREA 15.4081 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8334 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.69600425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.6299495 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 15.06 0.4 15.15 1.155 ;
    END
  END Q4N
  PIN D4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.66 0.625 11.805 0.905 ;
    END
  END D4
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1296 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 30 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.98 1.48 1.22 1.48 1.22 1.42 3.06 1.42 3.06 1.385 3.345 1.385 3.345 1.42 6.66 1.42 6.66 1.385 6.945 1.385 6.945 1.42 8.255 1.42 8.255 1.385 8.54 1.385 8.54 1.42 11.855 1.42 11.855 1.385 12.14 1.385 12.14 1.42 13.98 1.42 ;
    END
  END RN
  PIN Q3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.91405 LAYER Metal1 ;
    ANTENNADIFFAREA 13.53865 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8334 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.69600425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.6299495 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.95 0.765 10.91 0.765 10.91 1.18 10.85 1.18 10.85 0.4 10.95 0.4 ;
    END
  END Q3
  PIN Q3N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.91405 LAYER Metal1 ;
    ANTENNADIFFAREA 14.04855 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8334 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.69600425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.6299495 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.46 0.4 11.55 1.155 ;
    END
  END Q3N
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.06 0.625 8.205 0.905 ;
    END
  END D3
  PIN Q2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.91405 LAYER Metal1 ;
    ANTENNADIFFAREA 14.280525 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8334 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.69600425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.6299495 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.35 1.18 4.29 1.18 4.29 0.765 4.25 0.765 4.25 0.4 4.35 0.4 ;
    END
  END Q2
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.91405 LAYER Metal1 ;
    ANTENNADIFFAREA 13.450625 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8334 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.69600425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.6299495 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.65 0.4 3.74 1.155 ;
    END
  END Q2N
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.995 0.625 7.14 0.905 ;
    END
  END D2
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.91405 LAYER Metal1 ;
    ANTENNADIFFAREA 12.5281 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8334 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.69600425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.6299495 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.75 1.18 0.69 1.18 0.69 0.765 0.65 0.765 0.65 0.4 0.75 0.4 ;
    END
  END Q1
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.91405 LAYER Metal1 ;
    ANTENNADIFFAREA 12.940725 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8334 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.69600425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.6299495 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.05 0.4 0.14 1.155 ;
    END
  END Q1N
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.395 0.625 3.54 0.905 ;
    END
  END D1
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.645 0.77 7.825 0.92 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.2 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.54 0.395 1.54 0.395 1.65 0.855 1.65 0.855 1.54 0.975 1.54 0.975 1.65 1.42 1.65 1.42 1.54 1.54 1.54 1.54 1.65 2.125 1.65 2.125 1.54 2.245 1.54 2.245 1.65 2.52 1.65 2.52 1.54 2.645 1.54 2.645 1.65 3.435 1.65 3.435 1.54 3.555 1.54 3.555 1.65 3.875 1.65 3.875 1.54 3.995 1.54 3.995 1.65 4.455 1.65 4.455 1.54 4.575 1.54 4.575 1.65 5.02 1.65 5.02 1.54 5.14 1.54 5.14 1.65 5.725 1.65 5.725 1.54 5.845 1.54 5.845 1.65 6.12 1.65 6.12 1.54 6.245 1.54 6.245 1.65 7.035 1.65 7.035 1.54 7.155 1.54 7.155 1.65 7.53 1.65 7.53 1.54 7.65 1.54 7.65 1.65 8.045 1.65 8.045 1.54 8.165 1.54 8.165 1.65 8.955 1.65 8.955 1.54 9.08 1.54 9.08 1.65 9.355 1.65 9.355 1.54 9.475 1.54 9.475 1.65 10.06 1.65 10.06 1.54 10.18 1.54 10.18 1.65 10.625 1.65 10.625 1.54 10.745 1.54 10.745 1.65 11.205 1.65 11.205 1.54 11.325 1.54 11.325 1.65 11.645 1.65 11.645 1.54 11.765 1.54 11.765 1.65 12.555 1.65 12.555 1.54 12.68 1.54 12.68 1.65 12.955 1.65 12.955 1.54 13.075 1.54 13.075 1.65 13.66 1.65 13.66 1.54 13.78 1.54 13.78 1.65 14.225 1.65 14.225 1.54 14.345 1.54 14.345 1.65 14.805 1.65 14.805 1.54 14.925 1.54 14.925 1.65 15.2 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.2 0.06 14.9 0.06 14.9 0.17 14.78 0.17 14.78 0.06 14.375 0.06 14.375 0.17 14.255 0.17 14.255 0.06 13.855 0.06 13.855 0.17 13.72 0.17 13.72 0.06 13 0.06 13 0.17 12.88 0.17 12.88 0.06 11.77 0.06 11.77 0.17 11.65 0.17 11.65 0.165 11.645 0.165 11.645 0.06 11.3 0.06 11.3 0.17 11.18 0.17 11.18 0.06 10.775 0.06 10.775 0.17 10.655 0.17 10.655 0.06 10.255 0.06 10.255 0.17 10.12 0.17 10.12 0.06 9.4 0.06 9.4 0.17 9.28 0.17 9.28 0.06 8.17 0.06 8.17 0.17 8.05 0.17 8.05 0.165 8.045 0.165 8.045 0.06 7.65 0.06 7.65 0.17 7.525 0.17 7.525 0.06 7.155 0.06 7.155 0.165 7.15 0.165 7.15 0.17 7.03 0.17 7.03 0.06 5.92 0.06 5.92 0.17 5.8 0.17 5.8 0.06 5.08 0.06 5.08 0.17 4.945 0.17 4.945 0.06 4.545 0.06 4.545 0.17 4.425 0.17 4.425 0.06 4.02 0.06 4.02 0.17 3.9 0.17 3.9 0.06 3.555 0.06 3.555 0.165 3.55 0.165 3.55 0.17 3.43 0.17 3.43 0.06 2.32 0.06 2.32 0.17 2.2 0.17 2.2 0.06 1.48 0.06 1.48 0.17 1.345 0.17 1.345 0.06 0.945 0.06 0.945 0.17 0.825 0.17 0.825 0.06 0.42 0.06 0.42 0.17 0.3 0.17 0.3 0.06 0 0.06 0 -0.06 15.2 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 14.98 0.86 14.92 0.86 14.92 0.83 14.73 0.83 14.73 1.02 14.67 1.02 14.67 0.54 14.73 0.54 14.73 0.77 14.92 0.77 14.92 0.74 14.98 0.74 ;
      POLYGON 14.385 0.83 14.2 0.83 14.2 1.12 13.69 1.12 13.69 0.765 13.75 0.765 13.75 1.06 14.14 1.06 14.14 0.49 13.995 0.49 13.995 0.43 14.2 0.43 14.2 0.77 14.385 0.77 ;
      POLYGON 14.05 0.715 13.99 0.715 13.99 0.685 13.61 0.685 13.61 1.025 13.46 1.025 13.46 1.115 13.4 1.115 13.4 0.965 13.55 0.965 13.55 0.47 13.47 0.47 13.47 0.5 13.41 0.5 13.41 0.375 13.47 0.375 13.47 0.41 13.61 0.41 13.61 0.625 13.99 0.625 13.99 0.595 14.05 0.595 ;
      POLYGON 13.995 0.3 13.33 0.3 13.33 0.615 13.49 0.615 13.49 0.885 13.43 0.885 13.43 0.675 13.27 0.675 13.27 0.3 12.565 0.3 12.565 0.39 12.505 0.39 12.505 0.3 12.055 0.3 12.055 0.855 11.995 0.855 11.995 0.3 11.74 0.3 11.74 0.325 11.645 0.325 11.645 0.3 9.73 0.3 9.73 0.615 9.89 0.615 9.89 0.885 9.83 0.885 9.83 0.675 9.67 0.675 9.67 0.3 8.965 0.3 8.965 0.39 8.905 0.39 8.905 0.3 8.455 0.3 8.455 0.855 8.395 0.855 8.395 0.3 8.14 0.3 8.14 0.325 8.045 0.325 8.045 0.3 7.4 0.3 7.4 1.1 7.26 1.1 7.26 0.77 7.34 0.77 7.34 0.3 7.155 0.3 7.155 0.325 7.06 0.325 7.06 0.3 6.805 0.3 6.805 0.855 6.745 0.855 6.745 0.3 6.295 0.3 6.295 0.39 6.235 0.39 6.235 0.3 5.53 0.3 5.53 0.675 5.37 0.675 5.37 0.885 5.31 0.885 5.31 0.615 5.47 0.615 5.47 0.3 3.555 0.3 3.555 0.325 3.46 0.325 3.46 0.3 3.205 0.3 3.205 0.855 3.145 0.855 3.145 0.3 2.695 0.3 2.695 0.39 2.635 0.39 2.635 0.3 1.93 0.3 1.93 0.675 1.77 0.675 1.77 0.885 1.71 0.885 1.71 0.615 1.87 0.615 1.87 0.3 1.205 0.3 1.205 0.24 1.87 0.24 1.87 0.185 1.93 0.185 1.93 0.24 5.47 0.24 5.47 0.185 5.53 0.185 5.53 0.24 9.67 0.24 9.67 0.185 9.73 0.185 9.73 0.24 13.27 0.24 13.27 0.185 13.33 0.185 13.33 0.24 13.995 0.24 ;
      POLYGON 13.98 1.36 12.23 1.36 12.23 1.3 11.775 1.3 11.775 1.36 8.63 1.36 8.63 1.3 8.175 1.3 8.175 1.36 7.025 1.36 7.025 1.3 6.57 1.3 6.57 1.36 3.425 1.36 3.425 1.3 2.97 1.3 2.97 1.36 1.22 1.36 1.22 1.3 2.88 1.3 2.88 1.24 3.425 1.24 3.425 1.195 3.54 1.195 3.54 1.3 6.48 1.3 6.48 1.24 7.025 1.24 7.025 1.195 7.14 1.195 7.14 1.3 7.5 1.3 7.5 0.895 7.46 0.895 7.46 0.495 7.56 0.495 7.56 0.625 7.765 0.625 7.765 0.505 7.825 0.505 7.825 0.705 7.56 0.705 7.56 1.005 7.855 1.005 7.855 1.065 7.56 1.065 7.56 1.3 8.06 1.3 8.06 1.195 8.175 1.195 8.175 1.24 8.72 1.24 8.72 1.3 11.66 1.3 11.66 1.195 11.775 1.195 11.775 1.24 12.32 1.24 12.32 1.3 13.98 1.3 ;
      POLYGON 13.21 1.09 13.15 1.09 13.15 0.71 12.58 0.71 12.58 0.65 13.15 0.65 13.15 0.38 13.21 0.38 ;
      POLYGON 13.07 0.895 13.01 0.895 13.01 0.87 12.175 0.87 12.175 1.15 12.115 1.15 12.115 0.81 12.345 0.81 12.345 0.46 12.405 0.46 12.405 0.81 13.01 0.81 13.01 0.775 13.07 0.775 ;
      RECT 12.285 1.04 12.84 1.1 ;
      RECT 11.865 0.46 11.925 1.14 ;
      POLYGON 11.38 0.86 11.32 0.86 11.32 0.83 11.13 0.83 11.13 1.02 11.07 1.02 11.07 0.54 11.13 0.54 11.13 0.77 11.32 0.77 11.32 0.74 11.38 0.74 ;
      POLYGON 10.785 0.83 10.6 0.83 10.6 1.12 10.09 1.12 10.09 0.765 10.15 0.765 10.15 1.06 10.54 1.06 10.54 0.49 10.395 0.49 10.395 0.43 10.6 0.43 10.6 0.77 10.785 0.77 ;
      POLYGON 10.45 0.715 10.39 0.715 10.39 0.685 10.01 0.685 10.01 1.025 9.86 1.025 9.86 1.115 9.8 1.115 9.8 0.965 9.95 0.965 9.95 0.47 9.87 0.47 9.87 0.5 9.81 0.5 9.81 0.375 9.87 0.375 9.87 0.41 10.01 0.41 10.01 0.625 10.39 0.625 10.39 0.595 10.45 0.595 ;
      POLYGON 9.61 1.09 9.55 1.09 9.55 0.71 8.98 0.71 8.98 0.65 9.55 0.65 9.55 0.38 9.61 0.38 ;
      POLYGON 9.47 0.895 9.41 0.895 9.41 0.87 8.575 0.87 8.575 1.15 8.515 1.15 8.515 0.81 8.745 0.81 8.745 0.46 8.805 0.46 8.805 0.81 9.41 0.81 9.41 0.775 9.47 0.775 ;
      RECT 8.685 1.04 9.24 1.1 ;
      RECT 8.265 0.46 8.325 1.14 ;
      RECT 6.875 0.46 6.935 1.14 ;
      POLYGON 6.685 1.15 6.625 1.15 6.625 0.87 5.79 0.87 5.79 0.895 5.73 0.895 5.73 0.775 5.79 0.775 5.79 0.81 6.395 0.81 6.395 0.46 6.455 0.46 6.455 0.81 6.685 0.81 ;
      RECT 5.96 1.04 6.515 1.1 ;
      POLYGON 6.22 0.71 5.65 0.71 5.65 1.09 5.59 1.09 5.59 0.38 5.65 0.38 5.65 0.65 6.22 0.65 ;
      POLYGON 5.4 1.115 5.34 1.115 5.34 1.025 5.19 1.025 5.19 0.685 4.81 0.685 4.81 0.715 4.75 0.715 4.75 0.595 4.81 0.595 4.81 0.625 5.19 0.625 5.19 0.41 5.33 0.41 5.33 0.375 5.39 0.375 5.39 0.5 5.33 0.5 5.33 0.47 5.25 0.47 5.25 0.965 5.4 0.965 ;
      POLYGON 5.11 1.12 4.6 1.12 4.6 0.83 4.415 0.83 4.415 0.77 4.6 0.77 4.6 0.43 4.805 0.43 4.805 0.49 4.66 0.49 4.66 1.06 5.05 1.06 5.05 0.765 5.11 0.765 ;
      POLYGON 4.13 1.02 4.07 1.02 4.07 0.83 3.88 0.83 3.88 0.86 3.82 0.86 3.82 0.74 3.88 0.74 3.88 0.77 4.07 0.77 4.07 0.54 4.13 0.54 ;
      RECT 3.275 0.46 3.335 1.14 ;
      POLYGON 3.085 1.15 3.025 1.15 3.025 0.87 2.19 0.87 2.19 0.895 2.13 0.895 2.13 0.775 2.19 0.775 2.19 0.81 2.795 0.81 2.795 0.46 2.855 0.46 2.855 0.81 3.085 0.81 ;
      RECT 2.36 1.04 2.915 1.1 ;
      POLYGON 2.62 0.71 2.05 0.71 2.05 1.09 1.99 1.09 1.99 0.38 2.05 0.38 2.05 0.65 2.62 0.65 ;
      POLYGON 1.8 1.115 1.74 1.115 1.74 1.025 1.59 1.025 1.59 0.685 1.21 0.685 1.21 0.715 1.15 0.715 1.15 0.595 1.21 0.595 1.21 0.625 1.59 0.625 1.59 0.41 1.73 0.41 1.73 0.375 1.79 0.375 1.79 0.5 1.73 0.5 1.73 0.47 1.65 0.47 1.65 0.965 1.8 0.965 ;
      POLYGON 1.51 1.12 1 1.12 1 0.83 0.815 0.83 0.815 0.77 1 0.77 1 0.43 1.205 0.43 1.205 0.49 1.06 0.49 1.06 1.06 1.45 1.06 1.45 0.765 1.51 0.765 ;
      POLYGON 0.53 1.02 0.47 1.02 0.47 0.83 0.28 0.83 0.28 0.86 0.22 0.86 0.22 0.74 0.28 0.74 0.28 0.77 0.47 0.77 0.47 0.54 0.53 0.54 ;
  END
END DFF4RX1

MACRO DFF4RX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFF4RX2 0 0 ;
  SIZE 16.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q4N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.61845 LAYER Metal1 ;
    ANTENNADIFFAREA 16.104325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0953 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.78156675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 65.05341 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 16.46 0.4 16.55 1.18 ;
    END
  END Q4N
  PIN Q4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.61845 LAYER Metal1 ;
    ANTENNADIFFAREA 16.370975 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0953 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.78156675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 65.05341 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.75 0.755 15.71 0.755 15.71 1.18 15.65 1.18 15.65 0.4 15.75 0.4 ;
    END
  END Q4
  PIN D4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.86 0.625 13.005 0.905 ;
    END
  END D4
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 26.20952375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.18 1.48 1.62 1.48 1.62 1.42 3.46 1.42 3.46 1.385 3.745 1.385 3.745 1.42 7.46 1.42 7.46 1.385 7.745 1.385 7.745 1.42 9.055 1.42 9.055 1.385 9.34 1.385 9.34 1.42 13.055 1.42 13.055 1.385 13.34 1.385 13.34 1.42 15.18 1.42 ;
    END
  END RN
  PIN Q3N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.61845 LAYER Metal1 ;
    ANTENNADIFFAREA 15.779525 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0953 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.78156675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 65.05341 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.46 0.4 12.55 1.18 ;
    END
  END Q3N
  PIN Q3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.61845 LAYER Metal1 ;
    ANTENNADIFFAREA 16.046175 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0953 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.78156675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 65.05341 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.75 0.755 11.71 0.755 11.71 1.18 11.65 1.18 11.65 0.4 11.75 0.4 ;
    END
  END Q3
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.86 0.625 9.005 0.905 ;
    END
  END D3
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.61845 LAYER Metal1 ;
    ANTENNADIFFAREA 16.647025 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0953 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.78156675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 65.05341 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.25 0.4 4.34 1.18 ;
    END
  END Q2N
  PIN Q2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.61845 LAYER Metal1 ;
    ANTENNADIFFAREA 13.89135 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0953 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.78156675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 65.05341 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.15 1.18 5.09 1.18 5.09 0.755 5.05 0.755 5.05 0.4 5.15 0.4 ;
    END
  END Q2
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.795 0.625 7.94 0.905 ;
    END
  END D2
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.61845 LAYER Metal1 ;
    ANTENNADIFFAREA 16.569475 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0953 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.78156675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 65.05341 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 0.4 0.34 1.18 ;
    END
  END Q1N
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 9.61845 LAYER Metal1 ;
    ANTENNADIFFAREA 16.0163 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0953 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.78156675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 65.05341 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.15 1.18 1.09 1.18 1.09 0.755 1.05 0.755 1.05 0.4 1.15 0.4 ;
    END
  END Q1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.795 0.625 3.94 0.905 ;
    END
  END D1
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.445 0.77 8.625 0.92 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.8 1.77 0 1.77 0 1.65 0.055 1.65 0.055 1.54 0.175 1.54 0.175 1.65 0.475 1.65 0.475 1.54 0.595 1.54 0.595 1.65 0.82 1.65 0.82 1.54 0.94 1.54 0.94 1.65 1.255 1.65 1.255 1.54 1.375 1.54 1.375 1.65 1.82 1.65 1.82 1.54 1.94 1.54 1.94 1.65 2.525 1.65 2.525 1.54 2.645 1.54 2.645 1.65 2.92 1.65 2.92 1.54 3.045 1.54 3.045 1.65 3.835 1.65 3.835 1.54 3.955 1.54 3.955 1.65 4.055 1.65 4.055 1.54 4.175 1.54 4.175 1.65 4.475 1.65 4.475 1.54 4.595 1.54 4.595 1.65 4.82 1.65 4.82 1.54 4.94 1.54 4.94 1.65 5.255 1.65 5.255 1.54 5.375 1.54 5.375 1.65 5.82 1.65 5.82 1.54 5.94 1.54 5.94 1.65 6.525 1.65 6.525 1.54 6.645 1.54 6.645 1.65 6.92 1.65 6.92 1.54 7.045 1.54 7.045 1.65 7.835 1.65 7.835 1.54 7.955 1.54 7.955 1.65 8.33 1.65 8.33 1.54 8.45 1.54 8.45 1.65 8.845 1.65 8.845 1.54 8.965 1.54 8.965 1.65 9.755 1.65 9.755 1.54 9.88 1.54 9.88 1.65 10.155 1.65 10.155 1.54 10.275 1.54 10.275 1.65 10.86 1.65 10.86 1.54 10.98 1.54 10.98 1.65 11.425 1.65 11.425 1.54 11.545 1.54 11.545 1.65 11.86 1.65 11.86 1.54 11.98 1.54 11.98 1.65 12.205 1.65 12.205 1.54 12.325 1.54 12.325 1.65 12.625 1.65 12.625 1.54 12.745 1.54 12.745 1.65 12.845 1.65 12.845 1.54 12.965 1.54 12.965 1.65 13.755 1.65 13.755 1.54 13.88 1.54 13.88 1.65 14.155 1.65 14.155 1.54 14.275 1.54 14.275 1.65 14.86 1.65 14.86 1.54 14.98 1.54 14.98 1.65 15.425 1.65 15.425 1.54 15.545 1.54 15.545 1.65 15.86 1.65 15.86 1.54 15.98 1.54 15.98 1.65 16.205 1.65 16.205 1.54 16.325 1.54 16.325 1.65 16.625 1.65 16.625 1.54 16.745 1.54 16.745 1.65 16.8 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 16.8 0.06 16.745 0.06 16.745 0.17 16.625 0.17 16.625 0.06 16.3 0.06 16.3 0.17 16.18 0.17 16.18 0.06 15.945 0.06 15.945 0.17 15.825 0.17 15.825 0.06 15.575 0.06 15.575 0.17 15.455 0.17 15.455 0.06 15.055 0.06 15.055 0.17 14.935 0.17 14.935 0.165 14.92 0.165 14.92 0.06 14.2 0.06 14.2 0.17 14.08 0.17 14.08 0.06 12.97 0.06 12.97 0.17 12.845 0.17 12.845 0.06 12.745 0.06 12.745 0.17 12.625 0.17 12.625 0.06 12.3 0.06 12.3 0.17 12.18 0.17 12.18 0.06 11.945 0.06 11.945 0.17 11.825 0.17 11.825 0.06 11.575 0.06 11.575 0.17 11.455 0.17 11.455 0.06 11.055 0.06 11.055 0.17 10.935 0.17 10.935 0.165 10.92 0.165 10.92 0.06 10.2 0.06 10.2 0.17 10.08 0.17 10.08 0.06 8.97 0.06 8.97 0.17 8.845 0.17 8.845 0.06 8.45 0.06 8.45 0.17 8.325 0.17 8.325 0.06 7.955 0.06 7.955 0.17 7.83 0.17 7.83 0.06 6.72 0.06 6.72 0.17 6.6 0.17 6.6 0.06 5.88 0.06 5.88 0.165 5.865 0.165 5.865 0.17 5.745 0.17 5.745 0.06 5.345 0.06 5.345 0.17 5.225 0.17 5.225 0.06 4.975 0.06 4.975 0.17 4.855 0.17 4.855 0.06 4.62 0.06 4.62 0.17 4.5 0.17 4.5 0.06 4.175 0.06 4.175 0.17 4.055 0.17 4.055 0.06 3.955 0.06 3.955 0.17 3.83 0.17 3.83 0.06 2.72 0.06 2.72 0.17 2.6 0.17 2.6 0.06 1.88 0.06 1.88 0.165 1.865 0.165 1.865 0.17 1.745 0.17 1.745 0.06 1.345 0.06 1.345 0.17 1.225 0.17 1.225 0.06 0.975 0.06 0.975 0.17 0.855 0.17 0.855 0.06 0.62 0.06 0.62 0.17 0.5 0.17 0.5 0.06 0.175 0.06 0.175 0.17 0.055 0.17 0.055 0.06 0 0.06 0 -0.06 16.8 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 16.38 0.86 16.32 0.86 16.32 0.83 16.13 0.83 16.13 1.02 16.07 1.02 16.07 0.54 16.13 0.54 16.13 0.77 16.32 0.77 16.32 0.74 16.38 0.74 ;
      POLYGON 15.585 0.83 15.45 0.83 15.45 1.12 14.89 1.12 14.89 0.765 14.95 0.765 14.95 1.06 15.39 1.06 15.39 0.49 15.195 0.49 15.195 0.43 15.45 0.43 15.45 0.77 15.585 0.77 ;
      POLYGON 15.285 0.7 14.81 0.7 14.81 1.025 14.66 1.025 14.66 1.115 14.6 1.115 14.6 0.965 14.75 0.965 14.75 0.47 14.67 0.47 14.67 0.5 14.61 0.5 14.61 0.375 14.67 0.375 14.67 0.41 14.81 0.41 14.81 0.64 15.285 0.64 ;
      POLYGON 15.195 0.3 14.53 0.3 14.53 0.615 14.69 0.615 14.69 0.885 14.63 0.885 14.63 0.675 14.47 0.675 14.47 0.3 13.765 0.3 13.765 0.39 13.705 0.39 13.705 0.3 13.255 0.3 13.255 0.855 13.195 0.855 13.195 0.3 12.94 0.3 12.94 0.325 12.845 0.325 12.845 0.3 10.53 0.3 10.53 0.615 10.69 0.615 10.69 0.885 10.63 0.885 10.63 0.675 10.47 0.675 10.47 0.3 9.765 0.3 9.765 0.39 9.705 0.39 9.705 0.3 9.255 0.3 9.255 0.855 9.195 0.855 9.195 0.3 8.94 0.3 8.94 0.325 8.845 0.325 8.845 0.3 8.2 0.3 8.2 1.1 8.06 1.1 8.06 0.77 8.14 0.77 8.14 0.3 7.955 0.3 7.955 0.325 7.86 0.325 7.86 0.3 7.605 0.3 7.605 0.855 7.545 0.855 7.545 0.3 7.095 0.3 7.095 0.39 7.035 0.39 7.035 0.3 6.33 0.3 6.33 0.675 6.17 0.675 6.17 0.885 6.11 0.885 6.11 0.615 6.27 0.615 6.27 0.3 3.955 0.3 3.955 0.325 3.86 0.325 3.86 0.3 3.605 0.3 3.605 0.855 3.545 0.855 3.545 0.3 3.095 0.3 3.095 0.39 3.035 0.39 3.035 0.3 2.33 0.3 2.33 0.675 2.17 0.675 2.17 0.885 2.11 0.885 2.11 0.615 2.27 0.615 2.27 0.3 1.605 0.3 1.605 0.24 2.27 0.24 2.27 0.185 2.33 0.185 2.33 0.24 6.27 0.24 6.27 0.185 6.33 0.185 6.33 0.24 10.47 0.24 10.47 0.185 10.53 0.185 10.53 0.24 14.47 0.24 14.47 0.185 14.53 0.185 14.53 0.24 15.195 0.24 ;
      POLYGON 15.18 1.36 13.43 1.36 13.43 1.3 12.975 1.3 12.975 1.36 9.43 1.36 9.43 1.3 8.975 1.3 8.975 1.36 7.825 1.36 7.825 1.3 7.37 1.3 7.37 1.36 3.825 1.36 3.825 1.3 3.37 1.3 3.37 1.36 1.62 1.36 1.62 1.3 3.28 1.3 3.28 1.24 3.825 1.24 3.825 1.195 3.94 1.195 3.94 1.3 7.28 1.3 7.28 1.24 7.825 1.24 7.825 1.195 7.94 1.195 7.94 1.3 8.3 1.3 8.3 0.895 8.26 0.895 8.26 0.495 8.36 0.495 8.36 0.625 8.565 0.625 8.565 0.505 8.625 0.505 8.625 0.705 8.36 0.705 8.36 1.005 8.655 1.005 8.655 1.065 8.36 1.065 8.36 1.3 8.86 1.3 8.86 1.195 8.975 1.195 8.975 1.24 9.52 1.24 9.52 1.3 12.86 1.3 12.86 1.195 12.975 1.195 12.975 1.24 13.52 1.24 13.52 1.3 15.18 1.3 ;
      POLYGON 14.41 1.09 14.35 1.09 14.35 0.71 13.78 0.71 13.78 0.65 14.35 0.65 14.35 0.38 14.41 0.38 ;
      POLYGON 14.27 0.895 14.21 0.895 14.21 0.87 13.375 0.87 13.375 1.15 13.315 1.15 13.315 0.81 13.545 0.81 13.545 0.46 13.605 0.46 13.605 0.81 14.21 0.81 14.21 0.775 14.27 0.775 ;
      RECT 13.485 1.04 14.04 1.1 ;
      RECT 13.065 0.46 13.125 1.14 ;
      POLYGON 12.38 0.86 12.32 0.86 12.32 0.83 12.13 0.83 12.13 1.02 12.07 1.02 12.07 0.54 12.13 0.54 12.13 0.77 12.32 0.77 12.32 0.74 12.38 0.74 ;
      POLYGON 11.585 0.83 11.45 0.83 11.45 1.12 10.89 1.12 10.89 0.765 10.95 0.765 10.95 1.06 11.39 1.06 11.39 0.49 11.195 0.49 11.195 0.43 11.45 0.43 11.45 0.77 11.585 0.77 ;
      POLYGON 11.285 0.7 10.81 0.7 10.81 1.025 10.66 1.025 10.66 1.115 10.6 1.115 10.6 0.965 10.75 0.965 10.75 0.47 10.67 0.47 10.67 0.5 10.61 0.5 10.61 0.375 10.67 0.375 10.67 0.41 10.81 0.41 10.81 0.64 11.285 0.64 ;
      POLYGON 10.41 1.09 10.35 1.09 10.35 0.71 9.78 0.71 9.78 0.65 10.35 0.65 10.35 0.38 10.41 0.38 ;
      POLYGON 10.27 0.895 10.21 0.895 10.21 0.87 9.375 0.87 9.375 1.15 9.315 1.15 9.315 0.81 9.545 0.81 9.545 0.46 9.605 0.46 9.605 0.81 10.21 0.81 10.21 0.775 10.27 0.775 ;
      RECT 9.485 1.04 10.04 1.1 ;
      RECT 9.065 0.46 9.125 1.14 ;
      RECT 7.675 0.46 7.735 1.14 ;
      POLYGON 7.485 1.15 7.425 1.15 7.425 0.87 6.59 0.87 6.59 0.895 6.53 0.895 6.53 0.775 6.59 0.775 6.59 0.81 7.195 0.81 7.195 0.46 7.255 0.46 7.255 0.81 7.485 0.81 ;
      RECT 6.76 1.04 7.315 1.1 ;
      POLYGON 7.02 0.71 6.45 0.71 6.45 1.09 6.39 1.09 6.39 0.38 6.45 0.38 6.45 0.65 7.02 0.65 ;
      POLYGON 6.2 1.115 6.14 1.115 6.14 1.025 5.99 1.025 5.99 0.7 5.515 0.7 5.515 0.64 5.99 0.64 5.99 0.41 6.13 0.41 6.13 0.375 6.19 0.375 6.19 0.5 6.13 0.5 6.13 0.47 6.05 0.47 6.05 0.965 6.2 0.965 ;
      POLYGON 5.91 1.12 5.35 1.12 5.35 0.83 5.215 0.83 5.215 0.77 5.35 0.77 5.35 0.43 5.605 0.43 5.605 0.49 5.41 0.49 5.41 1.06 5.85 1.06 5.85 0.765 5.91 0.765 ;
      POLYGON 4.73 1.02 4.67 1.02 4.67 0.83 4.48 0.83 4.48 0.86 4.42 0.86 4.42 0.74 4.48 0.74 4.48 0.77 4.67 0.77 4.67 0.54 4.73 0.54 ;
      RECT 3.675 0.46 3.735 1.14 ;
      POLYGON 3.485 1.15 3.425 1.15 3.425 0.87 2.59 0.87 2.59 0.895 2.53 0.895 2.53 0.775 2.59 0.775 2.59 0.81 3.195 0.81 3.195 0.46 3.255 0.46 3.255 0.81 3.485 0.81 ;
      RECT 2.76 1.04 3.315 1.1 ;
      POLYGON 3.02 0.71 2.45 0.71 2.45 1.09 2.39 1.09 2.39 0.38 2.45 0.38 2.45 0.65 3.02 0.65 ;
      POLYGON 2.2 1.115 2.14 1.115 2.14 1.025 1.99 1.025 1.99 0.7 1.515 0.7 1.515 0.64 1.99 0.64 1.99 0.41 2.13 0.41 2.13 0.375 2.19 0.375 2.19 0.5 2.13 0.5 2.13 0.47 2.05 0.47 2.05 0.965 2.2 0.965 ;
      POLYGON 1.91 1.12 1.35 1.12 1.35 0.83 1.215 0.83 1.215 0.77 1.35 0.77 1.35 0.43 1.605 0.43 1.605 0.49 1.41 0.49 1.41 1.06 1.85 1.06 1.85 0.765 1.91 0.765 ;
      POLYGON 0.73 1.02 0.67 1.02 0.67 0.83 0.48 0.83 0.48 0.86 0.42 0.86 0.42 0.74 0.48 0.74 0.48 0.77 0.67 0.77 0.67 0.54 0.73 0.54 ;
  END
END DFF4RX2

MACRO DFF4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFF4X1 0 0 ;
  SIZE 13.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.845 0.77 7.025 0.92 ;
    END
  END CK
  PIN Q2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.14215 LAYER Metal1 ;
    ANTENNADIFFAREA 11.4759 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8334 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.7697985 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 72.5053995 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.99 1.29 3.855 1.29 3.855 0.9 3.93 0.9 3.93 0.41 3.99 0.41 ;
    END
  END Q2
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.35185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.345 1.085 6.34 1.085 6.34 1.145 6.215 1.145 6.215 0.77 6.34 0.77 6.34 1.005 6.345 1.005 ;
    END
  END D2
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.14215 LAYER Metal1 ;
    ANTENNADIFFAREA 11.4759 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8334 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.7697985 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 72.5053995 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.35 1.29 3.29 1.29 3.29 0.93 3.26 0.93 3.26 0.6 3.29 0.6 3.29 0.41 3.35 0.41 ;
    END
  END Q2N
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.14215 LAYER Metal1 ;
    ANTENNADIFFAREA 10.5238 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8334 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.7697985 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 72.5053995 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.79 1.29 0.655 1.29 0.655 0.9 0.73 0.9 0.73 0.41 0.79 0.41 ;
    END
  END Q1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.25925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.015 0.77 3.14 1.145 ;
    END
  END D1
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.14215 LAYER Metal1 ;
    ANTENNADIFFAREA 10.5238 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8334 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.7697985 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 72.5053995 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.29 0.09 1.29 0.09 0.93 0.06 0.93 0.06 0.705 0.055 0.705 0.055 0.625 0.06 0.625 0.06 0.6 0.09 0.6 0.09 0.41 0.15 0.41 ;
    END
  END Q1N
  PIN Q4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.14215 LAYER Metal1 ;
    ANTENNADIFFAREA 10.5238 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8334 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.7697985 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 72.5053995 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.945 1.29 12.81 1.29 12.81 0.41 12.87 0.41 12.87 0.9 12.945 0.9 ;
    END
  END Q4
  PIN D4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.25925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.46 0.77 10.585 1.145 ;
    END
  END D4
  PIN Q4N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.14215 LAYER Metal1 ;
    ANTENNADIFFAREA 10.5238 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8334 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.7697985 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 72.5053995 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.54 0.93 13.51 0.93 13.51 1.29 13.45 1.29 13.45 0.41 13.51 0.41 13.51 0.6 13.54 0.6 ;
    END
  END Q4N
  PIN Q3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.14215 LAYER Metal1 ;
    ANTENNADIFFAREA 12.389375 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8334 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.7697985 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 72.5053995 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.745 1.29 9.61 1.29 9.61 0.41 9.67 0.41 9.67 0.9 9.745 0.9 ;
    END
  END Q3
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.25925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.26 0.77 7.385 1.145 ;
    END
  END D3
  PIN Q3N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.14215 LAYER Metal1 ;
    ANTENNADIFFAREA 12.389375 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8334 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.7697985 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 72.5053995 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.34 0.93 10.31 0.93 10.31 1.29 10.25 1.29 10.25 0.41 10.31 0.41 10.31 0.6 10.34 0.6 ;
    END
  END Q3N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.6 1.77 0 1.77 0 1.65 0.245 1.65 0.245 1.54 0.365 1.54 0.365 1.65 0.935 1.65 0.935 1.54 1.055 1.54 1.055 1.65 1.28 1.65 1.28 1.54 1.4 1.54 1.4 1.65 2.1 1.65 2.1 1.54 2.22 1.54 2.22 1.65 3.015 1.65 3.015 1.54 3.135 1.54 3.135 1.65 3.445 1.65 3.445 1.54 3.565 1.54 3.565 1.65 4.135 1.65 4.135 1.54 4.255 1.54 4.255 1.65 4.48 1.65 4.48 1.54 4.6 1.54 4.6 1.65 5.3 1.65 5.3 1.54 5.42 1.54 5.42 1.65 6.215 1.65 6.215 1.54 6.335 1.54 6.335 1.65 6.73 1.65 6.73 1.54 6.85 1.54 6.85 1.65 7.265 1.65 7.265 1.54 7.385 1.54 7.385 1.65 8.18 1.65 8.18 1.54 8.3 1.54 8.3 1.65 9 1.65 9 1.54 9.12 1.54 9.12 1.65 9.345 1.65 9.345 1.54 9.465 1.54 9.465 1.65 10.035 1.65 10.035 1.54 10.155 1.54 10.155 1.65 10.465 1.65 10.465 1.54 10.585 1.54 10.585 1.65 11.38 1.65 11.38 1.54 11.5 1.54 11.5 1.65 12.2 1.65 12.2 1.54 12.32 1.54 12.32 1.65 12.545 1.65 12.545 1.54 12.665 1.54 12.665 1.65 13.235 1.65 13.235 1.54 13.355 1.54 13.355 1.65 13.6 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.6 0.06 13.355 0.06 13.355 0.17 13.235 0.17 13.235 0.06 12.665 0.06 12.665 0.17 12.545 0.17 12.545 0.06 12.295 0.06 12.295 0.17 12.175 0.17 12.175 0.06 11.385 0.06 11.385 0.17 11.265 0.17 11.265 0.06 10.585 0.06 10.585 0.17 10.465 0.17 10.465 0.06 10.155 0.06 10.155 0.17 10.035 0.17 10.035 0.06 9.465 0.06 9.465 0.17 9.345 0.17 9.345 0.06 9.095 0.06 9.095 0.17 8.975 0.17 8.975 0.06 8.185 0.06 8.185 0.17 8.065 0.17 8.065 0.06 7.385 0.06 7.385 0.17 7.265 0.17 7.265 0.06 6.85 0.06 6.85 0.17 6.725 0.17 6.725 0.06 6.335 0.06 6.335 0.17 6.215 0.17 6.215 0.06 5.535 0.06 5.535 0.17 5.415 0.17 5.415 0.06 4.625 0.06 4.625 0.17 4.505 0.17 4.505 0.06 4.255 0.06 4.255 0.17 4.135 0.17 4.135 0.06 3.565 0.06 3.565 0.17 3.445 0.17 3.445 0.06 3.135 0.06 3.135 0.17 3.015 0.17 3.015 0.06 2.335 0.06 2.335 0.17 2.215 0.17 2.215 0.06 1.425 0.06 1.425 0.17 1.305 0.17 1.305 0.06 1.055 0.06 1.055 0.17 0.935 0.17 0.935 0.06 0.365 0.06 0.365 0.17 0.245 0.17 0.245 0.06 0 0.06 0 -0.06 13.6 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 13.37 0.82 13.31 0.82 13.31 0.79 13.09 0.79 13.09 1.02 13.03 1.02 13.03 0.54 13.09 0.54 13.09 0.7 13.37 0.7 ;
      POLYGON 12.71 0.82 12.65 0.82 12.65 0.68 12.47 0.68 12.47 1.21 12.41 1.21 12.41 0.765 12.225 0.765 12.225 0.825 12.165 0.825 12.165 0.705 12.41 0.705 12.41 0.47 12.47 0.47 12.47 0.62 12.71 0.62 ;
      POLYGON 12.345 0.985 12.105 0.985 12.105 1.18 11.835 1.18 11.835 1.12 12.045 1.12 12.045 0.6 11.845 0.6 11.845 0.54 12.105 0.54 12.105 0.925 12.285 0.925 12.285 0.865 12.345 0.865 ;
      POLYGON 12.09 0.31 11.775 0.31 11.775 0.79 11.945 0.79 11.945 1.035 11.885 1.035 11.885 0.85 11.715 0.85 11.715 0.31 11.08 0.31 11.08 0.44 11.02 0.44 11.02 0.345 10.78 0.345 10.78 0.31 8.575 0.31 8.575 0.79 8.745 0.79 8.745 1.035 8.685 1.035 8.685 0.85 8.515 0.85 8.515 0.31 7.88 0.31 7.88 0.44 7.82 0.44 7.82 0.345 7.58 0.345 7.58 0.31 6.6 0.31 6.6 1.1 6.46 1.1 6.46 0.77 6.54 0.77 6.54 0.31 6.02 0.31 6.02 0.345 5.78 0.345 5.78 0.44 5.72 0.44 5.72 0.31 5.085 0.31 5.085 0.85 4.915 0.85 4.915 1.035 4.855 1.035 4.855 0.79 5.025 0.79 5.025 0.31 2.82 0.31 2.82 0.345 2.58 0.345 2.58 0.44 2.52 0.44 2.52 0.31 1.885 0.31 1.885 0.85 1.715 0.85 1.715 1.035 1.655 1.035 1.655 0.79 1.825 0.79 1.825 0.31 1.51 0.31 1.51 0.25 2.52 0.25 2.52 0.22 2.82 0.22 2.82 0.25 5.72 0.25 5.72 0.22 6.02 0.22 6.02 0.25 7.58 0.25 7.58 0.22 7.88 0.22 7.88 0.25 10.78 0.25 10.78 0.22 11.08 0.22 11.08 0.25 12.09 0.25 ;
      POLYGON 11.945 1.48 1.655 1.48 1.655 1.42 1.825 1.42 1.825 0.93 1.885 0.93 1.885 1.42 2.665 1.42 2.665 0.695 2.725 0.695 2.725 1.385 3 1.385 3 1.42 5.025 1.42 5.025 0.93 5.085 0.93 5.085 1.42 5.865 1.42 5.865 0.695 5.925 0.695 5.925 1.385 6.2 1.385 6.2 1.42 6.66 1.42 6.66 0.495 6.76 0.495 6.76 0.625 6.965 0.625 6.965 0.505 7.025 0.505 7.025 0.705 6.76 0.705 6.76 1.005 7.055 1.005 7.055 1.065 6.74 1.065 6.74 1.42 7.4 1.42 7.4 1.385 7.675 1.385 7.675 0.695 7.735 0.695 7.735 1.42 8.515 1.42 8.515 0.93 8.575 0.93 8.575 1.42 10.6 1.42 10.6 1.385 10.875 1.385 10.875 0.695 10.935 0.695 10.935 1.42 11.715 1.42 11.715 0.93 11.775 0.93 11.775 1.42 11.945 1.42 ;
      POLYGON 11.655 1.22 11.595 1.22 11.595 0.785 11.305 0.785 11.305 0.725 11.59 0.725 11.59 0.475 11.655 0.475 ;
      POLYGON 11.48 1.005 11.42 1.005 11.42 0.945 11.235 0.945 11.235 1.18 11.035 1.18 11.035 1.12 11.175 1.12 11.175 0.63 10.955 0.63 10.955 0.51 11.015 0.51 11.015 0.57 11.235 0.57 11.235 0.885 11.48 0.885 ;
      RECT 10.73 0.48 10.79 1.22 ;
      POLYGON 10.17 0.82 10.11 0.82 10.11 0.79 9.89 0.79 9.89 1.02 9.83 1.02 9.83 0.54 9.89 0.54 9.89 0.7 10.17 0.7 ;
      POLYGON 9.51 0.82 9.45 0.82 9.45 0.68 9.27 0.68 9.27 1.21 9.21 1.21 9.21 0.765 9.025 0.765 9.025 0.825 8.965 0.825 8.965 0.705 9.21 0.705 9.21 0.47 9.27 0.47 9.27 0.62 9.51 0.62 ;
      POLYGON 9.145 0.985 8.905 0.985 8.905 1.18 8.635 1.18 8.635 1.12 8.845 1.12 8.845 0.6 8.645 0.6 8.645 0.54 8.905 0.54 8.905 0.925 9.085 0.925 9.085 0.865 9.145 0.865 ;
      POLYGON 8.455 1.22 8.395 1.22 8.395 0.785 8.105 0.785 8.105 0.725 8.39 0.725 8.39 0.475 8.455 0.475 ;
      POLYGON 8.28 1.005 8.22 1.005 8.22 0.945 8.035 0.945 8.035 1.18 7.835 1.18 7.835 1.12 7.975 1.12 7.975 0.63 7.755 0.63 7.755 0.51 7.815 0.51 7.815 0.57 8.035 0.57 8.035 0.885 8.28 0.885 ;
      RECT 7.53 0.48 7.59 1.22 ;
      RECT 6.01 0.48 6.07 1.22 ;
      POLYGON 5.845 0.63 5.625 0.63 5.625 1.12 5.765 1.12 5.765 1.18 5.565 1.18 5.565 0.945 5.38 0.945 5.38 1.005 5.32 1.005 5.32 0.885 5.565 0.885 5.565 0.57 5.785 0.57 5.785 0.51 5.845 0.51 ;
      POLYGON 5.495 0.785 5.205 0.785 5.205 1.22 5.145 1.22 5.145 0.475 5.21 0.475 5.21 0.725 5.495 0.725 ;
      POLYGON 4.965 1.18 4.695 1.18 4.695 0.985 4.455 0.985 4.455 0.865 4.515 0.865 4.515 0.925 4.695 0.925 4.695 0.54 4.955 0.54 4.955 0.6 4.755 0.6 4.755 1.12 4.965 1.12 ;
      POLYGON 4.635 0.825 4.575 0.825 4.575 0.765 4.39 0.765 4.39 1.21 4.33 1.21 4.33 0.68 4.15 0.68 4.15 0.82 4.09 0.82 4.09 0.62 4.33 0.62 4.33 0.47 4.39 0.47 4.39 0.705 4.635 0.705 ;
      POLYGON 3.77 1.02 3.71 1.02 3.71 0.79 3.49 0.79 3.49 0.82 3.43 0.82 3.43 0.7 3.71 0.7 3.71 0.54 3.77 0.54 ;
      RECT 2.81 0.48 2.87 1.22 ;
      POLYGON 2.645 0.63 2.425 0.63 2.425 1.12 2.565 1.12 2.565 1.18 2.365 1.18 2.365 0.945 2.18 0.945 2.18 1.005 2.12 1.005 2.12 0.885 2.365 0.885 2.365 0.57 2.585 0.57 2.585 0.51 2.645 0.51 ;
      POLYGON 2.295 0.785 2.005 0.785 2.005 1.22 1.945 1.22 1.945 0.475 2.01 0.475 2.01 0.725 2.295 0.725 ;
      POLYGON 1.765 1.18 1.495 1.18 1.495 0.985 1.255 0.985 1.255 0.865 1.315 0.865 1.315 0.925 1.495 0.925 1.495 0.54 1.755 0.54 1.755 0.6 1.555 0.6 1.555 1.12 1.765 1.12 ;
      POLYGON 1.435 0.825 1.375 0.825 1.375 0.765 1.19 0.765 1.19 1.21 1.13 1.21 1.13 0.68 0.95 0.68 0.95 0.82 0.89 0.82 0.89 0.62 1.13 0.62 1.13 0.47 1.19 0.47 1.19 0.705 1.435 0.705 ;
      POLYGON 0.57 1.02 0.51 1.02 0.51 0.79 0.29 0.79 0.29 0.82 0.23 0.82 0.23 0.7 0.51 0.7 0.51 0.54 0.57 0.54 ;
  END
END DFF4X1

MACRO DFF4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFF4X2 0 0 ;
  SIZE 15.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.645 0.77 7.825 0.92 ;
    END
  END CK
  PIN Q2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.99935 LAYER Metal1 ;
    ANTENNADIFFAREA 13.784925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0953 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.2163335 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 60.02738975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.66 4.64 0.66 4.64 0.9 4.8 0.9 4.8 1.29 4.74 1.29 4.74 1.085 4.58 1.085 4.58 0.595 4.74 0.595 4.74 0.41 4.8 0.41 ;
    END
  END Q2
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.25925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.015 0.77 7.14 1.145 ;
    END
  END D2
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.99935 LAYER Metal1 ;
    ANTENNADIFFAREA 13.784925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0953 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.2163335 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 60.02738975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.99 1.29 3.93 1.29 3.93 0.93 3.86 0.93 3.86 0.6 3.93 0.6 3.93 0.41 3.99 0.41 ;
    END
  END Q2N
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.99935 LAYER Metal1 ;
    ANTENNADIFFAREA 12.62965 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0953 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.2163335 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 60.02738975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.66 1.04 0.66 1.04 0.9 1.2 0.9 1.2 1.29 1.14 1.29 1.14 1.085 0.98 1.085 0.98 0.595 1.14 0.595 1.14 0.41 1.2 0.41 ;
    END
  END Q1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.25925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.415 0.77 3.54 1.145 ;
    END
  END D1
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.99935 LAYER Metal1 ;
    ANTENNADIFFAREA 12.62965 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0953 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.2163335 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 60.02738975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.39 1.29 0.33 1.29 0.33 0.93 0.26 0.93 0.26 0.705 0.255 0.705 0.255 0.625 0.26 0.625 0.26 0.6 0.33 0.6 0.33 0.41 0.39 0.41 ;
    END
  END Q1N
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.25925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.06 0.77 8.185 1.145 ;
    END
  END D3
  PIN Q3N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.99935 LAYER Metal1 ;
    ANTENNADIFFAREA 14.86915 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0953 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.2163335 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 60.02738975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.34 0.93 11.27 0.93 11.27 1.29 11.21 1.29 11.21 0.41 11.27 0.41 11.27 0.6 11.34 0.6 ;
    END
  END Q3N
  PIN Q3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.99935 LAYER Metal1 ;
    ANTENNADIFFAREA 14.86915 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0953 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.2163335 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 60.02738975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.62 1.085 10.46 1.085 10.46 1.29 10.4 1.29 10.4 0.9 10.56 0.9 10.56 0.66 10.4 0.66 10.4 0.41 10.46 0.41 10.46 0.595 10.62 0.595 ;
    END
  END Q3
  PIN D4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.35185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 11.785 1.145 11.66 1.145 11.66 1.085 11.655 1.085 11.655 1.005 11.66 1.005 11.66 0.77 11.785 0.77 ;
    END
  END D4
  PIN Q4N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.99935 LAYER Metal1 ;
    ANTENNADIFFAREA 12.62965 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0953 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.2163335 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 60.02738975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.94 0.93 14.87 0.93 14.87 1.29 14.81 1.29 14.81 0.41 14.87 0.41 14.87 0.6 14.94 0.6 ;
    END
  END Q4N
  PIN Q4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.99935 LAYER Metal1 ;
    ANTENNADIFFAREA 12.62965 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0953 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.2163335 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 60.02738975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 14.22 1.085 14.06 1.085 14.06 1.29 14 1.29 14 0.9 14.16 0.9 14.16 0.66 14 0.66 14 0.41 14.06 0.41 14.06 0.595 14.22 0.595 ;
    END
  END Q4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.2 1.77 0 1.77 0 1.65 0.115 1.65 0.115 1.54 0.235 1.54 0.235 1.65 0.485 1.65 0.485 1.54 0.605 1.54 0.605 1.65 0.94 1.65 0.94 1.54 1.06 1.54 1.06 1.65 1.28 1.65 1.28 1.54 1.4 1.54 1.4 1.65 1.735 1.65 1.735 1.54 1.855 1.54 1.855 1.65 2.5 1.65 2.5 1.54 2.62 1.54 2.62 1.65 3.415 1.65 3.415 1.54 3.535 1.54 3.535 1.65 3.715 1.65 3.715 1.54 3.835 1.54 3.835 1.65 4.085 1.65 4.085 1.54 4.205 1.54 4.205 1.65 4.54 1.65 4.54 1.54 4.66 1.54 4.66 1.65 4.88 1.65 4.88 1.54 5 1.54 5 1.65 5.335 1.65 5.335 1.54 5.455 1.54 5.455 1.65 6.1 1.65 6.1 1.54 6.22 1.54 6.22 1.65 7.015 1.65 7.015 1.54 7.135 1.54 7.135 1.65 7.53 1.65 7.53 1.54 7.65 1.54 7.65 1.65 8.065 1.65 8.065 1.54 8.185 1.54 8.185 1.65 8.98 1.65 8.98 1.54 9.1 1.54 9.1 1.65 9.745 1.65 9.745 1.54 9.865 1.54 9.865 1.65 10.2 1.65 10.2 1.54 10.32 1.54 10.32 1.65 10.54 1.65 10.54 1.54 10.66 1.54 10.66 1.65 10.995 1.65 10.995 1.54 11.115 1.54 11.115 1.65 11.365 1.65 11.365 1.54 11.485 1.54 11.485 1.65 11.665 1.65 11.665 1.54 11.785 1.54 11.785 1.65 12.58 1.65 12.58 1.54 12.7 1.54 12.7 1.65 13.345 1.65 13.345 1.54 13.465 1.54 13.465 1.65 13.8 1.65 13.8 1.54 13.92 1.54 13.92 1.65 14.14 1.65 14.14 1.54 14.26 1.54 14.26 1.65 14.595 1.65 14.595 1.54 14.715 1.54 14.715 1.65 14.965 1.65 14.965 1.54 15.085 1.54 15.085 1.65 15.2 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.2 0.06 15.085 0.06 15.085 0.17 14.965 0.17 14.965 0.06 14.715 0.06 14.715 0.17 14.595 0.17 14.595 0.06 14.26 0.06 14.26 0.17 14.14 0.17 14.14 0.06 13.92 0.06 13.92 0.17 13.8 0.17 13.8 0.06 13.495 0.06 13.495 0.17 13.375 0.17 13.375 0.06 12.585 0.06 12.585 0.17 12.465 0.17 12.465 0.06 11.785 0.06 11.785 0.17 11.665 0.17 11.665 0.06 11.485 0.06 11.485 0.17 11.365 0.17 11.365 0.06 11.115 0.06 11.115 0.17 10.995 0.17 10.995 0.06 10.66 0.06 10.66 0.17 10.54 0.17 10.54 0.06 10.32 0.06 10.32 0.17 10.2 0.17 10.2 0.06 9.895 0.06 9.895 0.17 9.775 0.17 9.775 0.06 8.985 0.06 8.985 0.17 8.865 0.17 8.865 0.06 8.185 0.06 8.185 0.17 8.065 0.17 8.065 0.06 7.65 0.06 7.65 0.17 7.525 0.17 7.525 0.06 7.135 0.06 7.135 0.17 7.015 0.17 7.015 0.06 6.335 0.06 6.335 0.17 6.215 0.17 6.215 0.06 5.425 0.06 5.425 0.17 5.305 0.17 5.305 0.06 5 0.06 5 0.17 4.88 0.17 4.88 0.06 4.66 0.06 4.66 0.17 4.54 0.17 4.54 0.06 4.205 0.06 4.205 0.17 4.085 0.17 4.085 0.06 3.835 0.06 3.835 0.17 3.715 0.17 3.715 0.06 3.535 0.06 3.535 0.17 3.415 0.17 3.415 0.06 2.735 0.06 2.735 0.17 2.615 0.17 2.615 0.06 1.825 0.06 1.825 0.17 1.705 0.17 1.705 0.06 1.4 0.06 1.4 0.17 1.28 0.17 1.28 0.06 1.06 0.06 1.06 0.17 0.94 0.17 0.94 0.06 0.605 0.06 0.605 0.17 0.485 0.17 0.485 0.06 0.235 0.06 0.235 0.17 0.115 0.17 0.115 0.06 0 0.06 0 -0.06 15.2 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 14.73 0.82 14.67 0.82 14.67 0.79 14.45 0.79 14.45 1.02 14.39 1.02 14.39 0.54 14.45 0.54 14.45 0.7 14.73 0.7 ;
      POLYGON 14.095 0.8 13.67 0.8 13.67 1.33 13.61 1.33 13.61 0.765 13.425 0.765 13.425 0.825 13.365 0.825 13.365 0.705 13.61 0.705 13.61 0.41 13.67 0.41 13.67 0.74 14.095 0.74 ;
      POLYGON 13.545 0.985 13.305 0.985 13.305 1.18 13.035 1.18 13.035 1.12 13.245 1.12 13.245 0.6 13.045 0.6 13.045 0.54 13.305 0.54 13.305 0.925 13.485 0.925 13.485 0.865 13.545 0.865 ;
      POLYGON 13.29 0.31 12.975 0.31 12.975 0.79 13.145 0.79 13.145 1.035 13.085 1.035 13.085 0.85 12.915 0.85 12.915 0.31 12.28 0.31 12.28 0.44 12.22 0.44 12.22 0.345 11.98 0.345 11.98 0.31 9.375 0.31 9.375 0.79 9.545 0.79 9.545 1.035 9.485 1.035 9.485 0.85 9.315 0.85 9.315 0.31 8.68 0.31 8.68 0.44 8.62 0.44 8.62 0.345 8.38 0.345 8.38 0.31 7.4 0.31 7.4 1.1 7.26 1.1 7.26 0.77 7.34 0.77 7.34 0.31 6.82 0.31 6.82 0.345 6.58 0.345 6.58 0.44 6.52 0.44 6.52 0.31 5.885 0.31 5.885 0.85 5.715 0.85 5.715 1.035 5.655 1.035 5.655 0.79 5.825 0.79 5.825 0.31 3.22 0.31 3.22 0.345 2.98 0.345 2.98 0.44 2.92 0.44 2.92 0.31 2.285 0.31 2.285 0.85 2.115 0.85 2.115 1.035 2.055 1.035 2.055 0.79 2.225 0.79 2.225 0.31 1.91 0.31 1.91 0.25 2.92 0.25 2.92 0.22 3.22 0.22 3.22 0.25 6.52 0.25 6.52 0.22 6.82 0.22 6.82 0.25 8.38 0.25 8.38 0.22 8.68 0.22 8.68 0.25 11.98 0.25 11.98 0.22 12.28 0.22 12.28 0.25 13.29 0.25 ;
      POLYGON 13.28 1.48 1.92 1.48 1.92 1.42 2.225 1.42 2.225 0.93 2.285 0.93 2.285 1.42 3.065 1.42 3.065 0.695 3.125 0.695 3.125 1.385 3.4 1.385 3.4 1.42 5.825 1.42 5.825 0.93 5.885 0.93 5.885 1.42 6.665 1.42 6.665 0.695 6.725 0.695 6.725 1.385 7 1.385 7 1.42 7.46 1.42 7.46 0.495 7.56 0.495 7.56 0.625 7.765 0.625 7.765 0.505 7.825 0.505 7.825 0.705 7.56 0.705 7.56 1.005 7.855 1.005 7.855 1.065 7.54 1.065 7.54 1.42 8.2 1.42 8.2 1.385 8.475 1.385 8.475 0.695 8.535 0.695 8.535 1.42 9.315 1.42 9.315 0.93 9.375 0.93 9.375 1.42 11.8 1.42 11.8 1.385 12.075 1.385 12.075 0.695 12.135 0.695 12.135 1.42 12.915 1.42 12.915 0.93 12.975 0.93 12.975 1.42 13.28 1.42 ;
      POLYGON 12.855 1.22 12.795 1.22 12.795 0.785 12.505 0.785 12.505 0.725 12.79 0.725 12.79 0.475 12.855 0.475 ;
      POLYGON 12.68 1.005 12.62 1.005 12.62 0.945 12.435 0.945 12.435 1.18 12.235 1.18 12.235 1.12 12.375 1.12 12.375 0.63 12.155 0.63 12.155 0.51 12.215 0.51 12.215 0.57 12.435 0.57 12.435 0.885 12.68 0.885 ;
      RECT 11.93 0.48 11.99 1.22 ;
      POLYGON 11.13 0.82 11.07 0.82 11.07 0.79 10.85 0.79 10.85 1.02 10.79 1.02 10.79 0.54 10.85 0.54 10.85 0.7 11.13 0.7 ;
      POLYGON 10.495 0.8 10.07 0.8 10.07 1.33 10.01 1.33 10.01 0.765 9.825 0.765 9.825 0.825 9.765 0.825 9.765 0.705 10.01 0.705 10.01 0.41 10.07 0.41 10.07 0.74 10.495 0.74 ;
      POLYGON 9.945 0.985 9.705 0.985 9.705 1.18 9.435 1.18 9.435 1.12 9.645 1.12 9.645 0.6 9.445 0.6 9.445 0.54 9.705 0.54 9.705 0.925 9.885 0.925 9.885 0.865 9.945 0.865 ;
      POLYGON 9.255 1.22 9.195 1.22 9.195 0.785 8.905 0.785 8.905 0.725 9.19 0.725 9.19 0.475 9.255 0.475 ;
      POLYGON 9.08 1.005 9.02 1.005 9.02 0.945 8.835 0.945 8.835 1.18 8.635 1.18 8.635 1.12 8.775 1.12 8.775 0.63 8.555 0.63 8.555 0.51 8.615 0.51 8.615 0.57 8.835 0.57 8.835 0.885 9.08 0.885 ;
      RECT 8.33 0.48 8.39 1.22 ;
      RECT 6.81 0.48 6.87 1.22 ;
      POLYGON 6.645 0.63 6.425 0.63 6.425 1.12 6.565 1.12 6.565 1.18 6.365 1.18 6.365 0.945 6.18 0.945 6.18 1.005 6.12 1.005 6.12 0.885 6.365 0.885 6.365 0.57 6.585 0.57 6.585 0.51 6.645 0.51 ;
      POLYGON 6.295 0.785 6.005 0.785 6.005 1.22 5.945 1.22 5.945 0.475 6.01 0.475 6.01 0.725 6.295 0.725 ;
      POLYGON 5.765 1.18 5.495 1.18 5.495 0.985 5.255 0.985 5.255 0.865 5.315 0.865 5.315 0.925 5.495 0.925 5.495 0.54 5.755 0.54 5.755 0.6 5.555 0.6 5.555 1.12 5.765 1.12 ;
      POLYGON 5.435 0.825 5.375 0.825 5.375 0.765 5.19 0.765 5.19 1.33 5.13 1.33 5.13 0.8 4.705 0.8 4.705 0.74 5.13 0.74 5.13 0.41 5.19 0.41 5.19 0.705 5.435 0.705 ;
      POLYGON 4.41 1.02 4.35 1.02 4.35 0.79 4.13 0.79 4.13 0.82 4.07 0.82 4.07 0.7 4.35 0.7 4.35 0.54 4.41 0.54 ;
      RECT 3.21 0.48 3.27 1.22 ;
      POLYGON 3.045 0.63 2.825 0.63 2.825 1.12 2.965 1.12 2.965 1.18 2.765 1.18 2.765 0.945 2.58 0.945 2.58 1.005 2.52 1.005 2.52 0.885 2.765 0.885 2.765 0.57 2.985 0.57 2.985 0.51 3.045 0.51 ;
      POLYGON 2.695 0.785 2.405 0.785 2.405 1.22 2.345 1.22 2.345 0.475 2.41 0.475 2.41 0.725 2.695 0.725 ;
      POLYGON 2.165 1.18 1.895 1.18 1.895 0.985 1.655 0.985 1.655 0.865 1.715 0.865 1.715 0.925 1.895 0.925 1.895 0.54 2.155 0.54 2.155 0.6 1.955 0.6 1.955 1.12 2.165 1.12 ;
      POLYGON 1.835 0.825 1.775 0.825 1.775 0.765 1.59 0.765 1.59 1.33 1.53 1.33 1.53 0.8 1.105 0.8 1.105 0.74 1.53 0.74 1.53 0.41 1.59 0.41 1.59 0.705 1.835 0.705 ;
      POLYGON 0.81 1.02 0.75 1.02 0.75 0.79 0.53 0.79 0.53 0.82 0.47 0.82 0.47 0.7 0.75 0.7 0.75 0.54 0.81 0.54 ;
  END
END DFF4X2

MACRO DFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQX1 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8768 LAYER Metal1 ;
    ANTENNADIFFAREA 2.055125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.23085 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.1299545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 64.39896025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.14 0.73 0.13 0.73 0.13 1.375 0.07 1.375 0.07 0.73 0.06 0.73 0.06 0.59 0.07 0.59 0.07 0.52 0.13 0.52 0.13 0.59 0.14 0.59 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.04854375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.57 0.735 2.8 0.895 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.29629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.475 1.11 0.235 1.11 0.235 0.98 0.395 0.98 0.395 0.74 0.475 0.74 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.255 0.335 1.255 0.335 1.65 0.895 1.65 0.895 1.315 1.015 1.315 1.015 1.65 1.84 1.65 1.84 1.325 1.965 1.325 1.965 1.65 2.655 1.65 2.655 1.03 2.715 1.03 2.715 1.65 3.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 0.06 2.775 0.06 2.775 0.315 2.655 0.315 2.655 0.06 1.935 0.06 1.935 0.29 1.875 0.29 1.875 0.06 1.01 0.06 1.01 0.41 0.95 0.41 0.95 0.06 0.335 0.06 0.335 0.5 0.275 0.5 0.275 0.06 0 0.06 0 -0.06 3.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.98 1.085 2.92 1.085 2.92 0.475 2.495 0.475 2.495 0.305 2.21 0.305 2.21 0.655 2.15 0.655 2.15 0.455 1.755 0.455 1.755 0.285 1.565 0.285 1.565 0.695 1.29 0.695 1.29 0.865 1.23 0.865 1.23 0.63 1.505 0.63 1.505 0.225 1.815 0.225 1.815 0.395 2.15 0.395 2.15 0.245 2.555 0.245 2.555 0.415 2.92 0.415 2.92 0.355 2.98 0.355 ;
      POLYGON 2.86 0.635 2.47 0.635 2.47 1.245 2.18 1.245 2.18 1.345 2.24 1.345 2.24 1.405 2.12 1.405 2.12 1.245 0.605 1.245 0.605 1.375 0.49 1.375 0.49 1.255 0.545 1.255 0.545 0.52 0.605 0.52 0.605 1.185 1.5 1.185 1.5 0.775 1.56 0.775 1.56 1.185 2.41 1.185 2.41 0.575 2.86 0.575 ;
      POLYGON 2.35 0.855 2.275 0.855 2.275 1.085 2.215 1.085 2.215 0.855 1.78 0.855 1.78 0.735 1.84 0.735 1.84 0.795 2.29 0.795 2.29 0.365 2.35 0.365 ;
      POLYGON 2.04 0.665 1.98 0.665 1.98 0.605 1.695 0.605 1.695 1.085 1.635 1.085 1.635 0.375 1.695 0.375 1.695 0.545 2.04 0.545 ;
      POLYGON 1.395 0.465 1.17 0.465 1.17 0.965 1.38 0.965 1.38 1.085 1.32 1.085 1.32 1.025 0.82 1.025 0.82 0.67 0.88 0.67 0.88 0.965 1.11 0.965 1.11 0.405 1.395 0.405 ;
      POLYGON 1.05 0.865 0.99 0.865 0.99 0.57 0.745 0.57 0.745 1.085 0.685 1.085 0.685 0.42 0.455 0.42 0.455 0.66 0.29 0.66 0.29 0.8 0.23 0.8 0.23 0.6 0.395 0.6 0.395 0.36 0.805 0.36 0.805 0.51 1.05 0.51 ;
  END
END DFFHQX1

MACRO DFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQX2 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1834 LAYER Metal1 ;
    ANTENNADIFFAREA 2.536725 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2601 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.39446375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 67.42791225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.375 0.98 3.34 0.98 3.34 1.465 3.28 1.465 3.28 1.11 3.26 1.11 3.26 0.98 3.28 0.98 3.28 0.92 3.315 0.92 3.315 0.54 3.375 0.54 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.045 0.885 0.965 0.885 0.965 1.085 0.745 1.085 0.745 0.805 1.045 0.805 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.285 0.895 0.205 0.895 0.205 0.73 0.06 0.73 0.06 0.54 0.14 0.54 0.14 0.65 0.285 0.65 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 0 1.77 0 1.65 0.18 1.65 0.18 0.995 0.24 0.995 0.24 1.65 0.81 1.65 0.81 1.345 0.87 1.345 0.87 1.65 1.88 1.65 1.88 1.54 2 1.54 2 1.65 3.075 1.65 3.075 1.21 3.135 1.21 3.135 1.65 3.485 1.65 3.485 1.08 3.545 1.08 3.545 1.65 4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.695 0.06 3.695 0.575 3.635 0.575 3.635 0.06 2.995 0.06 2.995 0.485 3.055 0.485 3.055 0.545 2.935 0.545 2.935 0.06 1.855 0.06 1.855 0.485 1.915 0.485 1.915 0.545 1.795 0.545 1.795 0.06 1.055 0.06 1.055 0.545 0.935 0.545 0.935 0.485 0.995 0.485 0.995 0.06 0.28 0.06 0.28 0.2 0.22 0.2 0.22 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.9 0.98 3.78 0.98 3.78 1.385 3.72 1.385 3.72 0.98 3.475 0.98 3.475 0.86 3.535 0.86 3.535 0.92 3.84 0.92 3.84 0.54 3.9 0.54 ;
      POLYGON 3.715 0.82 3.655 0.82 3.655 0.735 3.475 0.735 3.475 0.44 3.215 0.44 3.215 0.705 2.97 0.705 2.97 1.245 2.715 1.245 2.715 1.465 2.655 1.465 2.655 1.185 2.91 1.185 2.91 0.705 2.775 0.705 2.775 0.63 2.625 0.63 2.625 0.57 2.835 0.57 2.835 0.645 3.155 0.645 3.155 0.38 3.535 0.38 3.535 0.675 3.715 0.675 ;
      POLYGON 2.81 0.865 2.395 0.865 2.395 1.085 2.335 1.085 2.335 0.44 2.075 0.44 2.075 0.705 1.695 0.705 1.695 1.055 1.635 1.055 1.635 0.47 1.215 0.47 1.215 0.95 1.145 0.95 1.145 0.705 0.775 0.705 0.775 0.47 0.445 0.47 0.445 1.02 0.385 1.02 0.385 0.41 0.715 0.41 0.715 0.385 0.835 0.385 0.835 0.645 1.155 0.645 1.155 0.41 1.695 0.41 1.695 0.645 2.015 0.645 2.015 0.38 2.395 0.38 2.395 0.805 2.81 0.805 ;
      POLYGON 2.65 1.085 2.555 1.085 2.555 1.435 1.315 1.435 1.315 1.245 0.665 1.245 0.665 1.37 0.555 1.37 0.555 0.57 0.675 0.57 0.675 0.63 0.615 0.63 0.615 1.185 1.315 1.185 1.315 0.985 1.375 0.985 1.375 1.375 2.495 1.375 2.495 1.025 2.59 1.025 2.59 0.965 2.65 0.965 ;
      POLYGON 2.295 1.245 2.175 1.245 2.175 0.865 1.795 0.865 1.795 0.805 2.175 0.805 2.175 0.54 2.235 0.54 2.235 1.185 2.295 1.185 ;
      POLYGON 2.075 1.215 1.535 1.215 1.535 1.275 1.475 1.275 1.475 0.63 1.315 0.63 1.315 0.57 1.535 0.57 1.535 1.155 2.015 1.155 2.015 0.965 2.075 0.965 ;
  END
END DFFHQX2

MACRO DFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQX4 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.1 0.815 4.6 0.895 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.43 0.34 0.93 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.70485 LAYER Metal1 ;
    ANTENNADIFFAREA 3.218175 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.341775 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.91412475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 62.96247525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.15 1.29 1.09 1.29 1.09 0.99 1.045 0.99 1.045 0.73 0.74 0.73 0.74 1.29 0.68 1.29 0.68 0.73 0.66 0.73 0.66 0.63 0.545 0.63 0.545 0.57 0.74 0.57 0.74 0.67 1.045 0.67 1.045 0.54 1.105 0.54 1.105 0.93 1.15 0.93 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.475 1.65 0.475 0.9 0.535 0.9 0.535 1.65 0.885 1.65 0.885 0.9 0.945 0.9 0.945 1.65 1.335 1.65 1.335 0.91 1.395 0.91 1.395 1.65 2.04 1.65 2.04 0.985 2.1 0.985 2.1 1.65 3.255 1.65 3.255 1.315 3.315 1.315 3.315 1.65 4.23 1.65 4.23 1.155 4.29 1.155 4.29 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 4.395 0.06 4.395 0.555 4.335 0.555 4.335 0.06 3.44 0.06 3.44 0.4 3.32 0.4 3.32 0.34 3.38 0.34 3.38 0.06 2.245 0.06 2.245 0.405 2.125 0.405 2.125 0.345 2.185 0.345 2.185 0.06 1.425 0.06 1.425 0.39 1.485 0.39 1.485 0.45 1.365 0.45 1.365 0.06 0.9 0.06 0.9 0.17 0.78 0.17 0.78 0.06 0.43 0.06 0.43 0.17 0.31 0.17 0.31 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.76 1.055 4 1.055 4 1.26 3.56 1.26 3.56 1.215 2.84 1.215 2.84 1.405 2.36 1.405 2.36 1.345 2.78 1.345 2.78 0.77 2.9 0.77 2.9 0.83 2.84 0.83 2.84 1.155 3.62 1.155 3.62 1.2 3.94 1.2 3.94 0.895 3.88 0.895 3.88 0.835 4 0.835 4 0.995 4.7 0.995 4.7 0.555 4.54 0.555 4.54 0.435 4.6 0.435 4.6 0.495 4.76 0.495 ;
      POLYGON 4.54 0.715 4.06 0.715 4.06 0.655 4.165 0.655 4.165 0.39 3.61 0.39 3.61 0.82 3.62 0.82 3.62 0.88 3.5 0.88 3.5 0.82 3.55 0.82 3.55 0.56 3.16 0.56 3.16 0.39 2.46 0.39 2.46 0.65 2.52 0.65 2.52 0.71 2.4 0.71 2.4 0.565 1.965 0.565 1.965 0.39 1.645 0.39 1.645 0.61 1.205 0.61 1.205 0.33 0.16 0.33 0.16 1.03 0.3 1.03 0.3 1.15 0.24 1.15 0.24 1.09 0.1 1.09 0.1 0.27 1.265 0.27 1.265 0.55 1.585 0.55 1.585 0.33 2.025 0.33 2.025 0.505 2.4 0.505 2.4 0.33 3.22 0.33 3.22 0.5 3.55 0.5 3.55 0.33 4.225 0.33 4.225 0.655 4.54 0.655 ;
      POLYGON 4.065 0.55 3.78 0.55 3.78 1.1 3.72 1.1 3.72 1.04 3.34 1.04 3.34 0.895 3.16 0.895 3.16 0.835 3.4 0.835 3.4 0.98 3.72 0.98 3.72 0.49 4.065 0.49 ;
      POLYGON 3.45 0.72 3.06 0.72 3.06 1.055 2.94 1.055 2.94 0.995 3 0.995 3 0.55 2.94 0.55 2.94 0.49 3.06 0.49 3.06 0.66 3.45 0.66 ;
      POLYGON 2.68 0.885 2.515 0.885 2.515 1.245 2.455 1.245 2.455 0.885 1.935 0.885 1.935 0.825 2.62 0.825 2.62 0.55 2.56 0.55 2.56 0.49 2.68 0.49 ;
      POLYGON 2.3 0.725 1.835 0.725 1.835 1.275 1.775 1.275 1.775 0.77 1.265 0.77 1.265 0.83 1.205 0.83 1.205 0.71 1.745 0.71 1.745 0.49 1.865 0.49 1.865 0.55 1.805 0.55 1.805 0.665 2.3 0.665 ;
  END
END DFFHQX4

MACRO DFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQX8 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.77777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.04 0.67 5.19 0.94 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.94 0.94 4.86 0.94 4.86 0.92 4.63 0.92 4.63 0.67 4.71 0.67 4.71 0.785 4.94 0.785 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.0392 LAYER Metal1 ;
    ANTENNADIFFAREA 3.738925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.499275 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.0872265 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 48.27399725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.37 1.345 1.31 1.345 1.31 0.66 0.96 0.66 0.96 1.345 0.9 1.345 0.9 0.66 0.55 0.66 0.55 1.345 0.49 1.345 0.49 0.73 0.14 0.73 0.14 1.345 0.08 1.345 0.08 0.73 0.06 0.73 0.06 0.6 0.08 0.6 0.08 0.54 0.14 0.54 0.14 0.67 0.49 0.67 0.49 0.54 0.55 0.54 0.55 0.6 0.9 0.6 0.9 0.54 0.96 0.54 0.96 0.6 1.31 0.6 1.31 0.54 1.37 0.54 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 1.77 0 1.77 0 1.65 0.285 1.65 0.285 0.9 0.345 0.9 0.345 1.65 0.695 1.65 0.695 0.9 0.755 0.9 0.755 1.65 1.105 1.65 1.105 0.9 1.165 0.9 1.165 1.65 1.515 1.65 1.515 0.955 1.575 0.955 1.575 1.65 1.925 1.65 1.925 1.33 2.045 1.33 2.045 1.39 1.985 1.39 1.985 1.65 2.615 1.65 2.615 1.54 2.735 1.54 2.735 1.65 3.83 1.65 3.83 1.365 3.95 1.365 3.95 1.425 3.89 1.425 3.89 1.65 4.57 1.65 4.57 1.2 4.69 1.2 4.69 1.26 4.63 1.26 4.63 1.65 5.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 0.06 4.765 0.06 4.765 0.41 4.705 0.41 4.705 0.06 3.89 0.06 3.89 0.285 3.95 0.285 3.95 0.345 3.83 0.345 3.83 0.06 2.75 0.06 2.75 0.32 2.81 0.32 2.81 0.38 2.69 0.38 2.69 0.06 1.985 0.06 1.985 0.52 1.925 0.52 1.925 0.06 1.575 0.06 1.575 0.52 1.515 0.52 1.515 0.06 1.165 0.06 1.165 0.485 1.105 0.485 1.105 0.06 0.755 0.06 0.755 0.485 0.695 0.485 0.695 0.06 0.345 0.06 0.345 0.485 0.285 0.485 0.285 0.06 0 0.06 0 -0.06 5.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.23 0.435 4.925 0.435 4.925 0.57 4.53 0.57 4.53 1.04 5.175 1.04 5.175 1.16 5.115 1.16 5.115 1.1 4.43 1.1 4.43 1.42 4.05 1.42 4.05 1.265 3.51 1.265 3.51 1.39 2.455 1.39 2.455 1.33 3.45 1.33 3.45 0.765 3.51 0.765 3.51 1.205 4.11 1.205 4.11 1.36 4.37 1.36 4.37 1.04 4.47 1.04 4.47 0.51 4.865 0.51 4.865 0.375 5.17 0.375 5.17 0.315 5.23 0.315 ;
      POLYGON 4.37 0.9 4.27 0.9 4.27 1.26 4.21 1.26 4.21 0.9 3.77 0.9 3.77 0.84 4.31 0.84 4.31 0.375 4.37 0.375 ;
      POLYGON 4.21 0.665 4.15 0.665 4.15 0.505 3.67 0.505 3.67 0.305 3.35 0.305 3.35 0.725 3.28 0.725 3.28 0.605 3.29 0.605 3.29 0.305 2.97 0.305 2.97 0.915 2.5 0.915 2.5 1.07 2.38 1.07 2.38 1.01 2.44 1.01 2.44 0.855 2.91 0.855 2.91 0.54 2.485 0.54 2.485 0.375 2.545 0.375 2.545 0.48 2.91 0.48 2.91 0.245 3.73 0.245 3.73 0.445 4.21 0.445 ;
      POLYGON 4.05 0.665 3.67 0.665 3.67 1.105 3.61 1.105 3.61 0.665 3.45 0.665 3.45 0.405 3.57 0.405 3.57 0.605 4.05 0.605 ;
      POLYGON 3.19 0.465 3.13 0.465 3.13 1.23 2 1.23 2 0.86 1.94 0.86 1.94 0.8 2.06 0.8 2.06 1.17 3.07 1.17 3.07 0.405 3.19 0.405 ;
      POLYGON 2.81 0.7 2.22 0.7 2.22 0.985 2.28 0.985 2.28 1.045 2.16 1.045 2.16 0.7 1.78 0.7 1.78 1.345 1.72 1.345 1.72 0.76 1.53 0.76 1.53 0.82 1.47 0.82 1.47 0.7 1.72 0.7 1.72 0.54 1.78 0.54 1.78 0.64 2.13 0.64 2.13 0.54 2.19 0.54 2.19 0.64 2.81 0.64 ;
  END
END DFFHQX8

MACRO DFFNSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRX1 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.173875 LAYER Metal1 ;
    ANTENNADIFFAREA 3.1741 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2529 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.549921 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 99.51364175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.765 1.11 0.74 1.11 0.74 1.345 0.68 1.345 0.68 1.11 0.635 1.11 0.635 0.45 0.68 0.45 0.68 0.41 0.74 0.41 0.74 0.53 0.695 0.53 0.695 0.955 0.765 0.955 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.173875 LAYER Metal1 ;
    ANTENNADIFFAREA 3.1741 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2529 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.549921 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 99.51364175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.14 0.54 0.13 0.54 0.13 1.29 0.05 1.29 0.05 0.405 0.14 0.405 ;
    END
  END QN
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.962963 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.17 0.92 5.155 0.92 5.155 0.99 5.075 0.99 5.075 0.92 5.025 0.92 5.025 0.79 5.075 0.79 5.075 0.705 5.155 0.705 5.155 0.79 5.17 0.79 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.9444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.595 0.815 4.58 0.815 4.58 0.945 4.5 0.945 4.5 0.73 4.435 0.73 4.435 0.6 4.5 0.6 4.5 0.46 4.595 0.46 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 25.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.62 1.495 3.56 1.495 3.56 1.325 3.215 1.325 3.215 1.23 1.665 1.23 1.665 0.93 1.66 0.93 1.66 0.73 1.74 0.73 1.74 0.93 1.725 0.93 1.725 1.17 3.275 1.17 3.275 1.265 3.62 1.265 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.81481475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.025 1.125 0.945 1.125 0.945 0.92 0.835 0.92 0.835 0.785 1.025 0.785 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 1.77 0 1.77 0 1.65 0.275 1.65 0.275 0.995 0.335 0.995 0.335 1.65 0.885 1.65 0.885 1.225 0.945 1.225 0.945 1.65 1.53 1.65 1.53 1.54 1.65 1.54 1.65 1.65 2.145 1.65 2.145 1.49 2.265 1.49 2.265 1.55 2.205 1.55 2.205 1.65 2.985 1.65 2.985 1.54 3.105 1.54 3.105 1.65 3.72 1.65 3.72 1.51 3.78 1.51 3.78 1.65 4.51 1.65 4.51 1.205 4.57 1.205 4.57 1.65 5.15 1.65 5.15 1.12 5.21 1.12 5.21 1.65 5.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 0.06 5.21 0.06 5.21 0.605 5.15 0.605 5.15 0.06 4.57 0.06 4.57 0.2 4.51 0.2 4.51 0.06 3.81 0.06 3.81 0.17 3.69 0.17 3.69 0.06 1.65 0.06 1.65 0.17 1.53 0.17 1.53 0.06 0.945 0.06 0.945 0.53 0.885 0.53 0.885 0.06 0.335 0.06 0.335 0.635 0.275 0.635 0.275 0.06 0 0.06 0 -0.06 5.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.005 0.72 4.945 0.72 4.945 1.025 5.005 1.025 5.005 1.425 4.945 1.425 4.945 1.085 4.885 1.085 4.885 0.66 4.945 0.66 4.945 0.36 3.54 0.36 3.54 0.305 2.855 0.305 2.855 0.245 3.6 0.245 3.6 0.3 5.005 0.3 ;
      POLYGON 4.835 0.6 4.775 0.6 4.775 1.23 4.715 1.23 4.715 1.105 4.37 1.105 4.37 1.36 3.745 1.36 3.745 1.205 3.335 1.205 3.335 1.085 3.015 1.085 3.015 0.835 3.075 0.835 3.075 1.025 3.395 1.025 3.395 1.145 3.805 1.145 3.805 1.3 4.31 1.3 4.31 0.925 4.105 0.925 4.105 0.985 4.045 0.985 4.045 0.865 4.31 0.865 4.31 0.81 4.37 0.81 4.37 1.045 4.715 1.045 4.715 0.54 4.835 0.54 ;
      POLYGON 4.27 0.6 3.985 0.6 3.985 1.14 4.175 1.14 4.175 1.2 3.925 1.2 3.925 0.765 3.39 0.765 3.39 0.705 3.925 0.705 3.925 0.54 4.27 0.54 ;
      POLYGON 3.865 0.925 3.515 0.925 3.515 1.025 3.575 1.025 3.575 1.085 3.455 1.085 3.455 0.925 3.255 0.925 3.255 0.73 2.94 0.73 2.94 1.05 2.795 1.05 2.795 0.99 2.88 0.99 2.88 0.73 2.855 0.73 2.855 0.49 2.915 0.49 2.915 0.67 3.26 0.67 3.26 0.485 3.32 0.485 3.32 0.865 3.865 0.865 ;
      POLYGON 3.575 0.575 3.42 0.575 3.42 0.425 3.115 0.425 3.115 0.605 3.055 0.605 3.055 0.365 3.48 0.365 3.48 0.515 3.575 0.515 ;
      POLYGON 3.285 1.465 3.095 1.465 3.095 1.39 2.045 1.39 2.045 1.45 1.985 1.45 1.985 1.39 1.125 1.39 1.125 0.435 1.185 0.435 1.185 1.33 3.155 1.33 3.155 1.405 3.285 1.405 ;
      POLYGON 2.82 0.9 2.735 0.9 2.735 0.395 2.525 0.395 2.525 0.335 2.795 0.335 2.795 0.78 2.82 0.78 ;
      POLYGON 2.675 1.08 2.615 1.08 2.615 0.89 1.8 0.89 1.8 0.65 1.515 0.65 1.515 0.855 1.455 0.855 1.455 0.59 1.86 0.59 1.86 0.83 2.615 0.83 2.615 0.49 2.675 0.49 ;
      RECT 1.785 0.99 2.5 1.05 ;
      POLYGON 2.47 0.71 2.005 0.71 2.005 0.455 2.07 0.455 2.07 0.65 2.41 0.65 2.41 0.49 2.47 0.49 ;
      POLYGON 2.27 0.55 2.21 0.55 2.21 0.395 1.905 0.395 1.905 0.52 1.77 0.52 1.77 0.46 1.845 0.46 1.845 0.335 2.27 0.335 ;
      POLYGON 1.955 0.275 1.75 0.275 1.75 0.335 1.385 0.335 1.385 1.05 1.325 1.05 1.325 0.31 1.065 0.31 1.065 0.685 0.755 0.685 0.755 0.625 1.005 0.625 1.005 0.25 1.69 0.25 1.69 0.215 1.955 0.215 ;
      POLYGON 0.54 1.02 0.46 1.02 0.46 0.815 0.19 0.815 0.19 0.735 0.46 0.735 0.46 0.54 0.54 0.54 ;
  END
END DFFNSRX1

MACRO DFFNSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRX2 0 0 ;
  SIZE 7 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.061625 LAYER Metal1 ;
    ANTENNADIFFAREA 4.01955 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318375 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.7573615 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 101.041225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.54 1.11 6.46 1.11 6.46 1.06 6.355 1.06 6.355 0.54 6.435 0.54 6.435 0.98 6.54 0.98 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.016025 LAYER Metal1 ;
    ANTENNADIFFAREA 4.01955 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318375 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.61413425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 100.42873975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.86 0.54 5.94 1.11 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 1.26 0.46 1.26 0.46 0.78 0.54 0.78 0.54 0.98 0.56 0.98 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.14 0.96 3.06 0.96 3.06 0.92 2.945 0.92 2.945 0.575 3.025 0.575 3.025 0.73 3.14 0.73 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.845 0.895 2.585 0.895 2.585 0.575 2.665 0.575 2.665 0.815 2.845 0.815 ;
    END
  END SN
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.36 1.26 0.28 1.26 0.28 0.92 0.26 0.92 0.26 0.78 0.34 0.78 0.34 0.79 0.36 0.79 ;
    END
  END CKN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7 1.77 0 1.77 0 1.65 0.36 1.65 0.36 1.36 0.42 1.36 0.42 1.65 1.34 1.65 1.34 1.51 1.4 1.51 1.4 1.65 1.725 1.65 1.725 1.51 1.785 1.51 1.785 1.65 2.54 1.65 2.54 1.54 2.66 1.54 2.66 1.65 4.425 1.65 4.425 1.235 4.485 1.235 4.485 1.65 4.79 1.65 4.79 1.2 4.94 1.2 4.94 1.14 5 1.14 5 1.26 4.85 1.26 4.85 1.65 5.54 1.65 5.54 1.355 5.6 1.355 5.6 1.65 6.225 1.65 6.225 1.51 6.285 1.51 6.285 1.65 6.695 1.65 6.695 1.51 6.755 1.51 6.755 1.65 7 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7 0.06 6.64 0.06 6.64 0.52 6.58 0.52 6.58 0.06 6.165 0.06 6.165 0.52 6.105 0.52 6.105 0.06 5.685 0.06 5.685 0.575 5.625 0.575 5.625 0.06 4.37 0.06 4.37 0.475 4.31 0.475 4.31 0.06 2.805 0.06 2.805 0.255 2.865 0.255 2.865 0.315 2.745 0.315 2.745 0.06 1.48 0.06 1.48 0.17 1.36 0.17 1.36 0.06 0.475 0.06 0.475 0.52 0.415 0.52 0.415 0.06 0 0.06 0 -0.06 7 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.92 1.07 6.86 1.07 6.86 0.68 6.595 0.68 6.595 0.83 6.535 0.83 6.535 0.62 6.83 0.62 6.83 0.425 6.89 0.425 6.89 0.62 6.92 0.62 ;
      POLYGON 6.76 1.27 5.7 1.27 5.7 1.255 5.365 1.255 5.365 1.465 4.95 1.465 4.95 1.405 5.305 1.405 5.305 1.195 5.7 1.195 5.7 0.735 5.42 0.735 5.42 0.54 5.48 0.54 5.48 0.675 5.76 0.675 5.76 1.21 6.04 1.21 6.04 0.72 6.1 0.72 6.1 1.21 6.7 1.21 6.7 0.78 6.76 0.78 ;
      POLYGON 5.44 0.955 3.85 0.955 3.85 1.13 3.79 1.13 3.79 0.54 3.85 0.54 3.85 0.895 5.38 0.895 5.38 0.835 5.44 0.835 ;
      POLYGON 5.11 0.635 4.63 0.635 4.63 0.39 4.71 0.39 4.71 0.555 5.03 0.555 5.03 0.39 5.11 0.39 ;
      POLYGON 4.965 0.795 3.95 0.795 3.95 0.315 3.08 0.315 3.08 0.415 3.3 0.415 3.3 0.93 3.36 0.93 3.36 0.99 3.24 0.99 3.24 0.475 2.585 0.475 2.585 0.22 2.395 0.22 2.395 0.16 2.645 0.16 2.645 0.415 3.02 0.415 3.02 0.255 4.01 0.255 4.01 0.735 4.965 0.735 ;
      POLYGON 4.93 0.455 4.81 0.455 4.81 0.29 4.53 0.29 4.53 0.635 4.11 0.635 4.11 0.515 4.17 0.515 4.17 0.575 4.47 0.575 4.47 0.23 4.87 0.23 4.87 0.395 4.93 0.395 ;
      POLYGON 4.69 1.26 4.61 1.26 4.61 1.135 3.965 1.135 3.965 1.055 4.69 1.055 ;
      POLYGON 3.945 1.415 3.825 1.415 3.825 1.31 2.92 1.31 2.92 1.28 2.265 1.28 2.265 0.88 1.7 0.88 1.7 0.82 2.325 0.82 2.325 1.22 2.98 1.22 2.98 1.25 3.63 1.25 3.63 0.72 3.69 0.72 3.69 1.25 3.885 1.25 3.885 1.355 3.945 1.355 ;
      POLYGON 3.725 1.47 2.76 1.47 2.76 1.44 2.105 1.44 2.105 1.115 1.505 1.115 1.505 0.98 0.98 0.98 0.98 0.92 1.54 0.92 1.54 0.66 1.505 0.66 1.505 0.54 1.565 0.54 1.565 0.6 1.6 0.6 1.6 1.055 2.165 1.055 2.165 1.38 2.82 1.38 2.82 1.41 3.725 1.41 ;
      POLYGON 3.53 1.15 3.08 1.15 3.08 1.12 2.425 1.12 2.425 0.635 1.71 0.635 1.71 0.33 1.14 0.33 1.14 0.27 1.77 0.27 1.77 0.575 2.075 0.575 2.075 0.38 2.135 0.38 2.135 0.575 2.485 0.575 2.485 1.025 2.545 1.025 2.545 1.06 3.14 1.06 3.14 1.09 3.47 1.09 3.47 0.54 3.53 0.54 ;
      POLYGON 2.37 0.445 2.235 0.445 2.235 0.28 1.93 0.28 1.93 0.475 1.87 0.475 1.87 0.22 2.295 0.22 2.295 0.385 2.37 0.385 ;
      POLYGON 2.005 1.375 0.88 1.375 0.88 1.385 0.82 1.385 0.82 0.425 0.88 0.425 0.88 1.315 2.005 1.315 ;
      POLYGON 1.44 0.805 0.98 0.805 0.98 0.325 0.72 0.325 0.72 1.115 0.66 1.115 0.66 0.68 0.16 0.68 0.16 1.265 0.18 1.265 0.18 1.385 0.12 1.385 0.12 1.315 0.1 1.315 0.1 0.46 0.21 0.46 0.21 0.4 0.27 0.4 0.27 0.52 0.16 0.52 0.16 0.62 0.66 0.62 0.66 0.265 1.04 0.265 1.04 0.745 1.44 0.745 ;
  END
END DFFNSRX2

MACRO DFFNSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRX4 0 0 ;
  SIZE 7.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.605575 LAYER Metal1 ;
    ANTENNADIFFAREA 4.788575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4716 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.76585025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 76.73028 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.185 0.565 6.655 0.565 6.655 0.86 6.95 0.86 6.95 1.33 6.89 1.33 6.89 0.92 6.54 0.92 6.54 1.33 6.48 1.33 6.48 0.92 6.26 0.92 6.26 0.79 6.34 0.79 6.34 0.86 6.595 0.86 6.595 0.505 7.185 0.505 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.605575 LAYER Metal1 ;
    ANTENNADIFFAREA 4.788575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4716 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.76585025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 76.73028 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.245 0.565 5.775 0.565 5.775 1.005 6.13 1.005 6.13 1.33 6.07 1.33 6.07 1.065 5.765 1.065 5.765 1.085 5.695 1.085 5.695 1.33 5.635 1.33 5.635 1.005 5.715 1.005 5.715 0.565 5.655 0.565 5.655 0.505 6.245 0.505 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.12 0.71 2.965 0.71 2.965 0.895 2.805 0.895 2.805 0.815 2.885 0.815 2.885 0.63 3.12 0.63 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.695 0.745 2.235 0.745 2.235 0.625 2.365 0.625 2.365 0.665 2.695 0.665 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.76 0.54 1.26 ;
    END
  END D
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.76 0.34 1.26 ;
    END
  END CKN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.8 1.77 0 1.77 0 1.65 0.395 1.65 0.395 1.36 0.455 1.36 0.455 1.65 1.25 1.65 1.25 1.51 1.31 1.51 1.31 1.65 1.825 1.65 1.825 1.54 1.945 1.54 1.945 1.65 2.46 1.65 2.46 1.54 2.58 1.54 2.58 1.65 4.425 1.65 4.425 1.24 4.545 1.24 4.545 1.3 4.485 1.3 4.485 1.65 4.97 1.65 4.97 1.21 5.03 1.21 5.03 1.65 5.405 1.65 5.405 1.02 5.465 1.02 5.465 1.65 5.865 1.65 5.865 1.165 5.925 1.165 5.925 1.65 6.275 1.65 6.275 1.145 6.335 1.145 6.335 1.65 6.685 1.65 6.685 1.02 6.745 1.02 6.745 1.65 7.12 1.65 7.12 1.01 7.18 1.01 7.18 1.65 7.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.8 0.06 7.505 0.06 7.505 0.455 7.445 0.455 7.445 0.06 6.95 0.06 6.95 0.17 6.83 0.17 6.83 0.06 6.48 0.06 6.48 0.17 6.36 0.17 6.36 0.06 6.01 0.06 6.01 0.17 5.89 0.17 5.89 0.06 5.395 0.06 5.395 0.51 5.335 0.51 5.335 0.06 4.985 0.06 4.985 0.51 4.925 0.51 4.925 0.06 3.075 0.06 3.075 0.37 2.955 0.37 2.955 0.31 3.015 0.31 3.015 0.06 1.46 0.06 1.46 0.17 1.34 0.17 1.34 0.06 0.455 0.06 0.455 0.5 0.395 0.5 0.395 0.06 0 0.06 0 -0.06 7.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.71 0.91 7.385 0.91 7.385 1.33 7.325 1.33 7.325 0.91 7.05 0.91 7.05 0.735 7.17 0.735 7.17 0.85 7.65 0.85 7.65 0.475 7.71 0.475 ;
      POLYGON 7.55 0.75 7.285 0.75 7.285 0.405 5.555 0.405 5.555 0.675 5.305 0.675 5.305 0.775 5.535 0.775 5.535 0.835 5.305 0.835 5.305 1.14 5.245 1.14 5.245 1.33 5.185 1.33 5.185 1.08 5.245 1.08 5.245 0.7 4.66 0.7 4.66 0.64 5.13 0.64 5.13 0.475 5.19 0.475 5.19 0.615 5.495 0.615 5.495 0.345 7.345 0.345 7.345 0.69 7.55 0.69 ;
      POLYGON 5.145 0.98 3.88 0.98 3.88 1.105 3.76 1.105 3.76 0.54 3.82 0.54 3.82 0.92 5.025 0.92 5.025 0.88 5.145 0.88 ;
      POLYGON 4.855 1.205 4.645 1.205 4.645 1.14 3.98 1.14 3.98 1.08 4.705 1.08 4.705 1.145 4.855 1.145 ;
      POLYGON 4.78 0.51 4.7 0.51 4.7 0.345 4.38 0.345 4.38 0.48 4.26 0.48 4.26 0.4 4.3 0.4 4.3 0.265 4.78 0.265 ;
      POLYGON 4.6 0.525 4.56 0.525 4.56 0.66 4 0.66 4 0.54 4.08 0.54 4.08 0.58 4.48 0.58 4.48 0.445 4.6 0.445 ;
      POLYGON 4.47 0.82 3.88 0.82 3.88 0.435 3.28 0.435 3.28 0.99 3.16 0.99 3.16 0.93 3.22 0.93 3.22 0.53 2.795 0.53 2.795 0.265 2.475 0.265 2.475 0.205 2.855 0.205 2.855 0.47 3.22 0.47 3.22 0.375 3.94 0.375 3.94 0.76 4.47 0.76 ;
      POLYGON 4 1.4 3.94 1.4 3.94 1.31 2.84 1.31 2.84 1.215 2.425 1.215 2.425 1.065 1.675 1.065 1.675 0.915 1.735 0.915 1.735 1.005 2.485 1.005 2.485 1.155 2.9 1.155 2.9 1.25 3.6 1.25 3.6 0.815 3.54 0.815 3.54 0.755 3.66 0.755 3.66 1.25 4 1.25 ;
      POLYGON 3.75 1.47 2.68 1.47 2.68 1.375 2.265 1.375 2.265 1.225 1.455 1.225 1.455 1.165 1.515 1.165 1.515 0.98 0.96 0.98 0.96 0.92 1.515 0.92 1.515 0.54 1.575 0.54 1.575 1.165 2.325 1.165 2.325 1.315 2.74 1.315 2.74 1.41 3.75 1.41 ;
      POLYGON 3.615 0.655 3.47 0.655 3.47 1.03 3.53 1.03 3.53 1.15 3 1.15 3 1.055 2.585 1.055 2.585 0.905 2.075 0.905 2.075 0.69 1.735 0.69 1.735 0.47 1.18 0.47 1.18 0.31 1.12 0.31 1.12 0.25 1.24 0.25 1.24 0.41 1.795 0.41 1.795 0.63 2.075 0.63 2.075 0.465 2.195 0.465 2.195 0.525 2.135 0.525 2.135 0.845 2.705 0.845 2.705 0.995 3.06 0.995 3.06 1.09 3.41 1.09 3.41 0.595 3.555 0.595 3.555 0.535 3.615 0.535 ;
      POLYGON 2.415 0.5 2.295 0.5 2.295 0.365 1.975 0.365 1.975 0.53 1.895 0.53 1.895 0.285 2.375 0.285 2.375 0.42 2.415 0.42 ;
      POLYGON 2.165 1.385 0.8 1.385 0.8 0.405 0.86 0.405 0.86 1.325 2.165 1.325 ;
      POLYGON 1.415 0.82 1.355 0.82 1.355 0.655 1.02 0.655 1.02 0.715 0.96 0.715 0.96 0.305 0.7 0.305 0.7 1.115 0.64 1.115 0.64 0.66 0.16 0.66 0.16 1.36 0.25 1.36 0.25 1.48 0.19 1.48 0.19 1.42 0.1 1.42 0.1 0.6 0.19 0.6 0.19 0.405 0.25 0.405 0.25 0.6 0.64 0.6 0.64 0.245 1.02 0.245 1.02 0.595 1.415 0.595 ;
  END
END DFFNSRX4

MACRO DFFNSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFNSRXL 0 0 ;
  SIZE 6.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.33165 LAYER Metal1 ;
    ANTENNADIFFAREA 3.350025 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2268 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.68981475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 112.9761905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.96 1.345 0.9 1.345 0.9 0.945 0.86 0.945 0.86 0.79 0.88 0.79 0.88 0.615 0.89 0.615 0.89 0.535 0.95 0.535 0.95 0.655 0.94 0.655 0.94 0.895 0.96 0.895 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.33165 LAYER Metal1 ;
    ANTENNADIFFAREA 3.350025 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2268 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.68981475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 112.9761905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.315 1.02 0.235 1.02 0.235 0.73 0.06 0.73 0.06 0.6 0.235 0.6 0.235 0.54 0.315 0.54 ;
    END
  END QN
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.17 0.895 6.09 0.895 6.09 0.705 5.915 0.705 5.915 0.57 6.17 0.57 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.39 0.975 5.31 0.975 5.31 0.73 5.25 0.73 5.25 0.535 5.33 0.535 5.33 0.6 5.39 0.6 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 29.212963 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.335 1.495 3.82 1.495 3.82 1.28 1.905 1.28 1.905 1.085 1.835 1.085 1.835 1.005 1.905 1.005 1.905 0.9 2.025 0.9 2.025 0.96 1.965 0.96 1.965 1.22 3.88 1.22 3.88 1.435 4.335 1.435 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.315 1.22 1.235 1.22 1.235 1.11 1.06 1.11 1.06 0.895 1.14 0.895 1.14 0.98 1.315 0.98 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 0 1.77 0 1.65 0.485 1.65 0.485 0.995 0.545 0.995 0.545 1.65 1.105 1.65 1.105 1.32 1.165 1.32 1.165 1.65 1.84 1.65 1.84 1.54 1.96 1.54 1.96 1.65 2.5 1.65 2.5 1.54 2.62 1.54 2.62 1.65 3.5 1.65 3.5 1.54 3.62 1.54 3.62 1.65 4.435 1.65 4.435 1.51 4.495 1.51 4.495 1.65 5.32 1.65 5.32 1.235 5.38 1.235 5.38 1.65 5.99 1.65 5.99 0.995 6.05 0.995 6.05 1.65 6.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 6.08 0.06 6.08 0.2 6.02 0.2 6.02 0.06 5.35 0.06 5.35 0.2 5.29 0.2 5.29 0.06 4.595 0.06 4.595 0.17 4.475 0.17 4.475 0.06 1.96 0.06 1.96 0.17 1.84 0.17 1.84 0.06 1.155 0.06 1.155 0.63 1.095 0.63 1.095 0.06 0.575 0.06 0.575 0.2 0.515 0.2 0.515 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.875 1.055 5.755 1.055 5.755 0.435 4.315 0.435 4.315 0.37 4.2 0.37 4.2 0.31 4.375 0.31 4.375 0.375 5.815 0.375 5.815 0.995 5.875 0.995 ;
      POLYGON 5.645 0.63 5.585 0.63 5.585 1.26 5.525 1.26 5.525 1.135 5.15 1.135 5.15 1.39 4.705 1.39 4.705 1.335 3.98 1.335 3.98 1.12 3.675 1.12 3.675 0.96 3.615 0.96 3.615 0.9 3.735 0.9 3.735 1.06 4.04 1.06 4.04 1.275 4.765 1.275 4.765 1.33 5.09 1.33 5.09 1.015 4.855 1.015 4.855 0.895 4.915 0.895 4.915 0.955 5.09 0.955 5.09 0.87 5.21 0.87 5.21 0.93 5.15 0.93 5.15 1.075 5.525 1.075 5.525 0.57 5.645 0.57 ;
      POLYGON 5.08 0.63 4.755 0.63 4.755 1.115 4.925 1.115 4.925 1.17 4.985 1.17 4.985 1.23 4.865 1.23 4.865 1.175 4.695 1.175 4.695 0.795 3.995 0.795 3.995 0.735 4.695 0.735 4.695 0.57 5.08 0.57 ;
      POLYGON 4.595 0.955 4.2 0.955 4.2 1.055 4.26 1.055 4.26 1.115 4.14 1.115 4.14 0.955 3.835 0.955 3.835 0.8 3.515 0.8 3.515 1.055 3.3 1.055 3.3 0.995 3.455 0.995 3.455 0.635 3.415 0.635 3.415 0.515 3.475 0.515 3.475 0.575 3.515 0.575 3.515 0.74 3.835 0.74 3.835 0.575 3.88 0.575 3.88 0.515 3.94 0.515 3.94 0.635 3.895 0.635 3.895 0.895 4.595 0.895 ;
      POLYGON 4.18 0.605 4.04 0.605 4.04 0.415 3.735 0.415 3.735 0.635 3.675 0.635 3.675 0.355 4.1 0.355 4.1 0.545 4.18 0.545 ;
      POLYGON 3.72 1.44 2.4 1.44 2.4 1.5 2.34 1.5 2.34 1.44 1.31 1.44 1.31 1.32 1.415 1.32 1.415 0.535 1.475 0.535 1.475 1.38 3.72 1.38 ;
      POLYGON 3.355 0.895 3.235 0.895 3.235 0.26 2.98 0.26 2.98 0.18 3.315 0.18 3.315 0.815 3.355 0.815 ;
      POLYGON 3.155 1.085 3.095 1.085 3.095 1.015 3.075 1.015 3.075 0.955 2.305 0.955 2.305 0.8 1.735 0.8 1.735 0.74 2.365 0.74 2.365 0.895 3.075 0.895 3.075 0.515 3.135 0.515 3.135 0.965 3.155 0.965 ;
      RECT 2.075 1.06 2.975 1.12 ;
      POLYGON 2.93 0.635 2.89 0.635 2.89 0.795 2.465 0.795 2.465 0.54 2.525 0.54 2.525 0.735 2.83 0.735 2.83 0.575 2.87 0.575 2.87 0.515 2.93 0.515 ;
      POLYGON 2.73 0.635 2.67 0.635 2.67 0.44 2.365 0.44 2.365 0.595 2.195 0.595 2.195 0.605 2.075 0.605 2.075 0.545 2.135 0.545 2.135 0.535 2.305 0.535 2.305 0.38 2.73 0.38 ;
      POLYGON 2.205 0.435 1.695 0.435 1.695 0.64 1.635 0.64 1.635 0.9 1.695 0.9 1.695 1.15 1.635 1.15 1.635 0.96 1.575 0.96 1.575 0.58 1.635 0.58 1.635 0.435 1.315 0.435 1.315 0.795 1.04 0.795 1.04 0.735 1.255 0.735 1.255 0.375 2.205 0.375 ;
      POLYGON 0.75 1.02 0.67 1.02 0.67 0.81 0.415 0.81 0.415 0.73 0.67 0.73 0.67 0.54 0.75 0.54 ;
  END
END DFFNSRXL

MACRO DFFQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFQX1 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.97105 LAYER Metal1 ;
    ANTENNADIFFAREA 1.93325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.17505 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.25992575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 89.04884325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.175 1.44 0.095 1.44 0.095 0.73 0.06 0.73 0.06 0.6 0.095 0.6 0.095 0.48 0.175 0.48 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.17 1.085 2.965 1.085 2.965 1.175 2.76 1.175 2.76 1.005 3.17 1.005 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.72 0.54 1.22 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 1.77 0 1.77 0 1.65 0.32 1.65 0.32 1.32 0.38 1.32 0.38 1.65 1.035 1.65 1.035 1.54 1.155 1.54 1.155 1.65 2.04 1.65 2.04 1.54 2.16 1.54 2.16 1.65 2.955 1.65 2.955 1.275 3.015 1.275 3.015 1.65 3.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 0.06 3.065 0.06 3.065 0.525 3.125 0.525 3.125 0.585 3.005 0.585 3.005 0.06 2.275 0.06 2.275 0.26 2.155 0.26 2.155 0.2 2.215 0.2 2.215 0.06 1.105 0.06 1.105 0.615 1.045 0.615 1.045 0.06 0.38 0.06 0.38 0.46 0.32 0.46 0.32 0.06 0 0.06 0 -0.06 3.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.33 1.3 3.27 1.3 3.27 0.745 2.845 0.745 2.845 0.42 1.735 0.42 1.735 0.85 1.81 0.85 1.81 0.91 1.495 0.91 1.495 1.08 1.435 1.08 1.435 0.85 1.675 0.85 1.675 0.36 2.905 0.36 2.905 0.685 3.24 0.685 3.24 0.52 3.3 0.52 3.3 0.685 3.33 0.685 ;
      POLYGON 3.17 0.905 2.66 0.905 2.66 1.43 1.655 1.43 1.655 1.46 1.255 1.46 1.255 1.44 0.59 1.44 0.59 1.32 0.64 1.32 0.64 0.48 0.7 0.48 0.7 1.38 1.315 1.38 1.315 1.4 1.595 1.4 1.595 1.05 1.715 1.05 1.715 1.11 1.655 1.11 1.655 1.37 2.6 1.37 2.6 1.085 2.4 1.085 2.4 0.965 2.46 0.965 2.46 1.025 2.6 1.025 2.6 0.845 2.675 0.845 2.675 0.785 2.735 0.785 2.735 0.845 3.17 0.845 ;
      POLYGON 2.695 0.685 2.3 0.685 2.3 1.21 2.5 1.21 2.5 1.27 2.24 1.27 2.24 0.96 2.13 0.96 2.13 1.02 2.07 1.02 2.07 0.9 2.24 0.9 2.24 0.625 2.635 0.625 2.635 0.52 2.695 0.52 ;
      POLYGON 2.14 0.8 1.97 0.8 1.97 1.27 1.805 1.27 1.805 1.21 1.91 1.21 1.91 0.75 1.835 0.75 1.835 0.52 1.895 0.52 1.895 0.69 1.97 0.69 1.97 0.74 2.08 0.74 2.08 0.68 2.14 0.68 ;
      POLYGON 1.575 0.61 1.335 0.61 1.335 1.18 1.495 1.18 1.495 1.3 1.435 1.3 1.435 1.24 1.275 1.24 1.275 1.07 1.02 1.07 1.02 1.01 1.275 1.01 1.275 0.55 1.575 0.55 ;
      POLYGON 1.175 0.91 0.92 0.91 0.92 1.27 0.8 1.27 0.8 1.21 0.84 1.21 0.84 0.38 0.54 0.38 0.54 0.62 0.335 0.62 0.335 0.76 0.275 0.76 0.275 0.56 0.48 0.56 0.48 0.32 0.9 0.32 0.9 0.85 1.175 0.85 ;
  END
END DFFQX1

MACRO DFFQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFQX2 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.07145 LAYER Metal1 ;
    ANTENNADIFFAREA 2.126825 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.211275 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.80452025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 78.714945 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.14 0.92 3.12 0.92 3.12 1.355 3.06 1.355 3.06 0.79 3.08 0.79 3.08 0.54 3.14 0.54 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.055 0.975 0.975 0.975 0.975 0.73 0.86 0.73 0.86 0.59 0.94 0.59 0.94 0.65 1.055 0.65 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.37 0.87 0.29 0.87 0.29 0.73 0.06 0.73 0.06 0.6 0.14 0.6 0.14 0.625 0.37 0.625 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 1.77 0 1.77 0 1.65 0.15 1.65 0.15 0.995 0.21 0.995 0.21 1.65 0.92 1.65 0.92 1.235 0.98 1.235 0.98 1.65 1.75 1.65 1.75 1.49 1.87 1.49 1.87 1.55 1.81 1.55 1.81 1.65 2.795 1.65 2.795 1.235 2.855 1.235 2.855 1.65 3.28 1.65 3.28 1.025 3.34 1.025 3.34 1.65 3.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 0.06 3.46 0.06 3.46 0.52 3.4 0.52 3.4 0.06 2.82 0.06 2.82 0.52 2.76 0.52 2.76 0.06 1.81 0.06 1.81 0.55 1.75 0.55 1.75 0.06 1.06 0.06 1.06 0.2 1 0.2 1 0.06 0.26 0.06 0.26 0.5 0.2 0.5 0.2 0.06 0 0.06 0 -0.06 3.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.665 0.925 3.545 0.925 3.545 1.275 3.485 1.275 3.485 0.925 3.24 0.925 3.24 0.805 3.3 0.805 3.3 0.865 3.605 0.865 3.605 0.485 3.665 0.485 ;
      POLYGON 3.505 0.765 3.445 0.765 3.445 0.705 3.24 0.705 3.24 0.44 2.98 0.44 2.98 0.68 2.45 0.68 2.45 1.17 2.51 1.17 2.51 1.23 2.39 1.23 2.39 0.485 2.51 0.485 2.51 0.62 2.92 0.62 2.92 0.38 3.3 0.38 3.3 0.645 3.505 0.645 ;
      POLYGON 2.67 1.39 1.155 1.39 1.155 1.135 0.775 1.135 0.775 1.26 0.7 1.26 0.7 0.52 0.64 0.52 0.64 0.43 0.76 0.43 0.76 1.075 1.155 1.075 1.155 0.97 1.215 0.97 1.215 1.33 2.61 1.33 2.61 1.07 2.55 1.07 2.55 0.95 2.61 0.95 2.61 1.01 2.67 1.01 ;
      POLYGON 2.585 0.35 2.29 0.35 2.29 0.985 2.23 0.985 2.23 0.355 1.97 0.355 1.97 0.71 1.595 0.71 1.595 1.07 1.475 1.07 1.475 1.01 1.535 1.01 1.535 0.36 0.84 0.36 0.84 0.33 0.53 0.33 0.53 1.02 0.47 1.02 0.47 0.27 0.9 0.27 0.9 0.3 1.24 0.3 1.24 0.24 1.36 0.24 1.36 0.3 1.595 0.3 1.595 0.65 1.91 0.65 1.91 0.295 2.255 0.295 2.255 0.29 2.585 0.29 ;
      POLYGON 2.25 1.23 2.07 1.23 2.07 0.87 1.695 0.87 1.695 0.81 2.07 0.81 2.07 0.455 2.13 0.455 2.13 1.17 2.25 1.17 ;
      POLYGON 1.955 1.23 1.315 1.23 1.315 0.485 1.435 0.485 1.435 0.545 1.375 0.545 1.375 1.17 1.895 1.17 1.895 0.97 1.955 0.97 ;
  END
END DFFQX2

MACRO DFFQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFQX4 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.765 0.895 3.565 0.895 3.565 0.975 3.485 0.975 3.485 0.675 3.565 0.675 3.565 0.815 3.765 0.815 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.46 0.34 0.96 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.32435 LAYER Metal1 ;
    ANTENNADIFFAREA 2.568175 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.29295 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.93428925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 62.140297 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.185 0.545 1.105 0.545 1.105 0.965 1.13 0.965 1.13 1.355 1.07 1.355 1.07 1.02 1.045 1.02 1.045 0.73 0.72 0.73 0.72 1.355 0.66 1.355 0.66 0.545 0.595 0.545 0.595 0.485 0.72 0.485 0.72 0.6 0.74 0.6 0.74 0.67 1.045 0.67 1.045 0.485 1.185 0.485 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 1.77 0 1.77 0 1.65 0.455 1.65 0.455 1.06 0.515 1.06 0.515 1.65 0.865 1.65 0.865 0.965 0.925 0.965 0.925 1.65 1.275 1.65 1.275 1.045 1.335 1.045 1.335 1.65 1.685 1.65 1.685 1.235 1.745 1.235 1.745 1.65 2.705 1.65 2.705 1.54 2.825 1.54 2.825 1.65 3.565 1.65 3.565 1.235 3.625 1.235 3.625 1.65 4.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 0.06 3.655 0.06 3.655 0.415 3.595 0.415 3.595 0.06 2.825 0.06 2.825 0.17 2.705 0.17 2.705 0.06 1.86 0.06 1.86 0.2 1.8 0.2 1.8 0.06 1.42 0.06 1.42 0.17 1.3 0.17 1.3 0.06 0.95 0.06 0.95 0.17 0.83 0.17 0.83 0.06 0.45 0.06 0.45 0.2 0.39 0.2 0.39 0.06 0 0.06 0 -0.06 4.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.005 0.545 3.945 0.545 3.945 0.875 3.925 0.875 3.925 1.26 3.77 1.26 3.77 1.135 3.38 1.135 3.38 1.39 2.31 1.39 2.31 1.065 2.12 1.065 2.12 0.945 2.18 0.945 2.18 1.005 2.385 1.005 2.385 0.805 2.445 0.805 2.445 1.065 2.37 1.065 2.37 1.33 3.32 1.33 3.32 0.98 3.38 0.98 3.38 1.075 3.865 1.075 3.865 0.815 3.885 0.815 3.885 0.485 4.005 0.485 ;
      POLYGON 3.785 0.715 3.665 0.715 3.665 0.575 3.385 0.575 3.385 0.745 3.325 0.745 3.325 0.355 3.06 0.355 3.06 0.98 3 0.98 3 0.355 2.115 0.355 2.115 0.36 0.16 0.36 0.16 1.06 0.31 1.06 0.31 1.18 0.25 1.18 0.25 1.12 0.1 1.12 0.1 0.3 2.055 0.3 2.055 0.295 3.385 0.295 3.385 0.515 3.725 0.515 3.725 0.655 3.785 0.655 ;
      POLYGON 3.22 1.23 2.84 1.23 2.84 1.06 2.705 1.06 2.705 1 2.9 1 2.9 1.17 3.16 1.17 3.16 0.455 3.22 0.455 ;
      POLYGON 2.9 0.77 2.605 0.77 2.605 1.23 2.47 1.23 2.47 1.17 2.545 1.17 2.545 0.545 2.47 0.545 2.47 0.485 2.605 0.485 2.605 0.71 2.84 0.71 2.84 0.65 2.9 0.65 ;
      POLYGON 2.285 0.845 2.02 0.845 2.02 1.17 2.2 1.17 2.2 1.23 1.96 1.23 1.96 0.995 1.64 0.995 1.64 0.875 1.7 0.875 1.7 0.935 1.96 0.935 1.96 0.785 2.225 0.785 2.225 0.455 2.285 0.455 ;
      POLYGON 1.86 0.835 1.8 0.835 1.8 0.775 1.54 0.775 1.54 1.355 1.48 1.355 1.48 0.775 1.205 0.775 1.205 0.715 1.595 0.715 1.595 0.545 1.535 0.545 1.535 0.485 1.655 0.485 1.655 0.715 1.86 0.715 ;
  END
END DFFQX4

MACRO DFFQXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFQXL 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8948 LAYER Metal1 ;
    ANTENNADIFFAREA 1.7432 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.69629625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 96.175926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.495 0.14 1.31 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.97 0.925 2.965 0.925 2.965 1.185 2.73 1.185 2.73 1.105 2.755 1.105 2.755 0.845 2.97 0.845 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.485 1.185 0.24 1.185 0.24 0.98 0.405 0.98 0.405 0.85 0.485 0.85 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.285 0.335 1.285 0.335 1.65 0.99 1.65 0.99 1.54 1.11 1.54 1.11 1.65 1.97 1.65 1.97 1.54 2.09 1.54 2.09 1.65 2.845 1.65 2.845 1.285 2.905 1.285 2.905 1.65 3.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 0.06 2.845 0.06 2.845 0.305 2.905 0.305 2.905 0.365 2.785 0.365 2.785 0.06 2.09 0.06 2.09 0.19 2.15 0.19 2.15 0.25 2.03 0.25 2.03 0.06 1.08 0.06 1.08 0.43 1.02 0.43 1.02 0.06 0.335 0.06 0.335 0.59 0.275 0.59 0.275 0.06 0 0.06 0 -0.06 3.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.13 1.31 3.07 1.31 3.07 0.525 2.625 0.525 2.625 0.235 2.31 0.235 2.31 0.41 1.87 0.41 1.87 0.235 1.61 0.235 1.61 0.67 1.745 0.67 1.745 0.73 1.44 0.73 1.44 1.085 1.38 1.085 1.38 0.67 1.55 0.67 1.55 0.175 1.93 0.175 1.93 0.35 2.25 0.35 2.25 0.175 2.685 0.175 2.685 0.465 3.05 0.465 3.05 0.335 3.13 0.335 ;
      POLYGON 2.97 0.745 2.63 0.745 2.63 1.44 1.62 1.44 1.62 1.47 1.24 1.47 1.24 1.44 0.585 1.44 0.585 0.85 0.595 0.85 0.595 0.495 0.655 0.495 0.655 0.89 0.645 0.89 0.645 1.38 1.3 1.38 1.3 1.41 1.56 1.41 1.56 1.03 1.62 1.03 1.62 1.38 2.57 1.38 2.57 1.055 2.33 1.055 2.33 0.935 2.39 0.935 2.39 0.995 2.57 0.995 2.57 0.685 2.605 0.685 2.605 0.625 2.665 0.625 2.665 0.685 2.97 0.685 ;
      POLYGON 2.525 0.455 2.47 0.455 2.47 0.8 2.23 0.8 2.23 1.22 2.47 1.22 2.47 1.28 2.17 1.28 2.17 0.8 2.065 0.8 2.065 0.86 2.005 0.86 2.005 0.74 2.41 0.74 2.41 0.395 2.465 0.395 2.465 0.335 2.525 0.335 ;
      POLYGON 2.07 0.64 1.905 0.64 1.905 1.28 1.735 1.28 1.735 1.22 1.845 1.22 1.845 0.57 1.71 0.57 1.71 0.335 1.77 0.335 1.77 0.51 1.905 0.51 1.905 0.58 2.01 0.58 2.01 0.52 2.07 0.52 ;
      POLYGON 1.46 1.31 1.4 1.31 1.4 1.245 1.22 1.245 1.22 0.87 0.975 0.87 0.975 0.75 1.035 0.75 1.035 0.81 1.22 0.81 1.22 0.365 1.45 0.365 1.45 0.425 1.28 0.425 1.28 1.185 1.46 1.185 ;
      POLYGON 1.12 0.65 0.875 0.65 0.875 1.28 0.755 1.28 0.755 1.22 0.815 1.22 0.815 0.395 0.495 0.395 0.495 0.75 0.3 0.75 0.3 0.81 0.24 0.81 0.24 0.69 0.435 0.69 0.435 0.335 0.875 0.335 0.875 0.59 1.06 0.59 1.06 0.53 1.12 0.53 ;
  END
END DFFQXL

MACRO DFFRHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRHQX1 0 0 ;
  SIZE 3.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.514725 LAYER Metal1 ;
    ANTENNADIFFAREA 2.20035 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.23085 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.893329 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 91.57894725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.14 1.16 0.13 1.16 0.13 1.36 0.065 1.36 0.065 1.16 0.06 1.16 0.06 0.425 0.065 0.425 0.065 0.28 0.13 0.28 0.13 0.555 0.12 0.555 0.12 0.905 0.13 0.905 0.13 0.965 0.14 0.965 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.7831715 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.08 0.79 1.365 0.935 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.79 0.455 0.92 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.76051775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.365 0.705 3.075 0.705 3.075 0.55 3.21 0.55 3.21 0.625 3.365 0.625 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1 0.335 1 0.335 1.65 0.72 1.65 0.72 1.12 0.78 1.12 0.78 1.65 1.2 1.65 1.2 1.155 1.26 1.155 1.26 1.65 2.065 1.65 2.065 1.15 2.125 1.15 2.125 1.65 2.475 1.65 2.475 1.12 2.535 1.12 2.535 1.65 3.235 1.65 3.235 1.14 3.295 1.14 3.295 1.65 3.6 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 0.06 3.305 0.06 3.305 0.305 3.365 0.305 3.365 0.365 3.235 0.365 3.235 0.06 3 0.06 3 0.305 3.06 0.305 3.06 0.365 2.94 0.365 2.94 0.06 2.125 0.06 2.125 0.425 2.065 0.425 2.065 0.06 1.24 0.06 1.24 0.43 1.18 0.43 1.18 0.06 0.335 0.06 0.335 0.52 0.275 0.52 0.275 0.06 0 0.06 0 -0.06 3.6 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.54 1.11 3.53 1.11 3.53 1.17 3.47 1.17 3.47 1.045 3.48 1.045 3.48 0.83 3.115 0.83 3.115 0.89 3.055 0.89 3.055 0.765 3.47 0.765 3.47 0.485 2.76 0.485 2.76 0.305 2.565 0.305 2.565 0.68 2.505 0.68 2.505 0.575 1.945 0.575 1.945 0.305 1.735 0.305 1.735 0.76 1.675 0.76 1.675 0.245 2.005 0.245 2.005 0.515 2.505 0.515 2.505 0.245 2.82 0.245 2.82 0.425 3.47 0.425 3.47 0.3 3.53 0.3 3.53 0.71 3.54 0.71 ;
      POLYGON 3.42 0.975 3.31 0.975 3.31 1.045 3.175 1.045 3.175 1.44 2.805 1.44 2.805 0.94 2.17 0.94 2.17 1.055 2.005 1.055 2.005 1.41 1.32 1.41 1.32 1.055 1.14 1.055 1.14 1.43 0.84 1.43 0.84 0.97 0.575 0.97 0.575 1.265 0.515 1.265 0.515 0.465 0.535 0.465 0.535 0.295 0.595 0.295 0.595 0.52 0.575 0.52 0.575 0.91 0.9 0.91 0.9 1.37 1.08 1.37 1.08 0.995 1.43 0.995 1.43 0.625 1.49 0.625 1.49 1.055 1.38 1.055 1.38 1.35 1.705 1.35 1.705 0.865 1.765 0.865 1.765 1.35 1.945 1.35 1.945 0.995 2.11 0.995 2.11 0.88 2.805 0.88 2.805 0.84 2.865 0.84 2.865 1.38 3.115 1.38 3.115 0.985 3.245 0.985 3.245 0.915 3.42 0.915 ;
      POLYGON 2.985 1.27 2.925 1.27 2.925 0.715 2.69 0.715 2.69 0.82 2.025 0.82 2.025 0.93 1.965 0.93 1.965 0.76 2.63 0.76 2.63 0.385 2.69 0.385 2.69 0.655 2.985 0.655 ;
      POLYGON 2.745 1.29 2.685 1.29 2.685 1.06 2.33 1.06 2.33 1.29 2.27 1.29 2.27 1 2.745 1 ;
      POLYGON 2.425 0.695 1.885 0.695 1.885 1.26 1.825 1.26 1.825 0.39 1.885 0.39 1.885 0.635 2.425 0.635 ;
      POLYGON 1.61 1.26 1.55 1.26 1.55 0.54 1.39 0.54 1.39 0.555 0.875 0.555 0.875 0.68 0.815 0.68 0.815 0.495 1.325 0.495 1.325 0.48 1.55 0.48 1.55 0.355 1.61 0.355 ;
      POLYGON 1.34 0.715 1.02 0.715 1.02 1.255 0.96 1.255 0.96 0.84 0.695 0.84 0.695 0.23 0.455 0.23 0.455 0.68 0.18 0.68 0.18 0.62 0.395 0.62 0.395 0.17 0.755 0.17 0.755 0.335 0.97 0.335 0.97 0.395 0.755 0.395 0.755 0.78 0.96 0.78 0.96 0.655 1.34 0.655 ;
  END
END DFFRHQX1

MACRO DFFRHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRHQX2 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6683 LAYER Metal1 ;
    ANTENNADIFFAREA 3.08665 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2601 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.25874675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 81.83391 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.53 0.34 1.305 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.75404525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.765 0.895 1.715 0.895 1.715 1.115 1.485 1.115 1.485 1.025 1.635 1.025 1.635 0.815 1.765 0.815 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.835 1.085 0.6 1.085 0.6 0.74 0.765 0.74 0.765 1.005 0.835 1.005 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.175 0.885 4.095 0.885 4.095 0.705 3.965 0.705 3.965 0.515 4.175 0.515 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.77 0 1.77 0 1.65 0.075 1.65 0.075 0.915 0.135 0.915 0.135 1.65 0.485 1.65 0.485 1.185 0.545 1.185 0.545 1.65 1.005 1.65 1.005 1.345 1.065 1.345 1.065 1.65 1.705 1.65 1.705 1.435 1.645 1.435 1.645 1.375 1.765 1.375 1.765 1.65 2.64 1.65 2.64 1.335 2.76 1.335 2.76 1.395 2.7 1.395 2.7 1.65 3.255 1.65 3.255 1.54 3.375 1.54 3.375 1.65 4.27 1.65 4.27 1.51 4.33 1.51 4.33 1.65 4.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 0.06 4.26 0.06 4.26 0.2 4.2 0.2 4.2 0.06 3.98 0.06 3.98 0.195 4.04 0.195 4.04 0.255 3.92 0.255 3.92 0.06 2.905 0.06 2.905 0.405 2.785 0.405 2.785 0.345 2.845 0.345 2.845 0.06 1.645 0.06 1.645 0.395 1.525 0.395 1.525 0.335 1.585 0.335 1.585 0.06 0.515 0.06 0.515 0.42 0.575 0.42 0.575 0.48 0.455 0.48 0.455 0.06 0.135 0.06 0.135 0.51 0.075 0.51 0.075 0.06 0 0.06 0 -0.06 4.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.5 1.325 4.44 1.325 4.44 1.265 4.17 1.265 4.17 1.425 2.86 1.425 2.86 1.235 2.305 1.235 2.305 1.28 1.865 1.28 1.865 1.275 1.545 1.275 1.545 1.435 1.165 1.435 1.165 1.245 0.755 1.245 0.755 1.305 0.695 1.305 0.695 1.185 0.935 1.185 0.935 0.415 0.995 0.415 0.995 1.185 1.225 1.185 1.225 1.375 1.485 1.375 1.485 1.215 1.865 1.215 1.865 0.715 1.805 0.715 1.805 0.655 1.925 0.655 1.925 1.22 2.245 1.22 2.245 0.9 2.185 0.9 2.185 0.84 2.305 0.84 2.305 1.175 2.92 1.175 2.92 1.365 3.645 1.365 3.645 1.045 3.585 1.045 3.585 0.985 3.705 0.985 3.705 1.365 4.11 1.365 4.11 1.205 4.5 1.205 ;
      POLYGON 4.495 1.105 4.435 1.105 4.435 1.045 3.965 1.045 3.965 0.985 4.275 0.985 4.275 0.415 3.76 0.415 3.76 0.405 3.44 0.405 3.44 0.665 3.5 0.665 3.5 0.725 3.38 0.725 3.38 0.565 2.625 0.565 2.625 0.405 2.245 0.405 2.245 0.665 2.305 0.665 2.305 0.725 2.185 0.725 2.185 0.345 2.685 0.345 2.685 0.505 3.38 0.505 3.38 0.345 3.82 0.345 3.82 0.355 4.335 0.355 4.335 0.985 4.435 0.985 4.435 0.54 4.495 0.54 ;
      POLYGON 3.865 1.235 3.805 1.235 3.805 0.885 2.74 0.885 2.74 0.945 2.68 0.945 2.68 0.825 3.6 0.825 3.6 0.565 3.54 0.565 3.54 0.505 3.66 0.505 3.66 0.825 3.865 0.825 ;
      POLYGON 3.545 1.265 3.02 1.265 3.02 1.185 3.465 1.185 3.465 1.145 3.545 1.145 ;
      POLYGON 3.28 0.725 2.525 0.725 2.525 1.075 2.405 1.075 2.405 1.015 2.465 1.015 2.465 0.565 2.405 0.565 2.405 0.505 2.525 0.505 2.525 0.665 3.28 0.665 ;
      POLYGON 2.145 1.12 2.085 1.12 2.085 1.06 2.025 1.06 2.025 0.555 1.375 0.555 1.375 0.64 1.255 0.64 1.255 0.58 1.315 0.58 1.315 0.495 2.025 0.495 2.025 0.39 2.085 0.39 2.085 1 2.145 1 ;
      POLYGON 1.705 0.715 1.535 0.715 1.535 0.8 1.385 0.8 1.385 1.275 1.325 1.275 1.325 0.8 1.095 0.8 1.095 0.415 1.155 0.415 1.155 0.315 0.835 0.315 0.835 0.64 0.5 0.64 0.5 0.82 0.44 0.82 0.44 0.58 0.775 0.58 0.775 0.255 1.215 0.255 1.215 0.475 1.155 0.475 1.155 0.74 1.475 0.74 1.475 0.655 1.705 0.655 ;
  END
END DFFRHQX2

MACRO DFFRHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRHQX4 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.069525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 16.3322545 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.74 0.85 3.3 0.85 3.3 0.365 2.415 0.365 2.415 0.555 2.095 0.555 2.095 0.715 2.035 0.715 2.035 0.555 1.94 0.555 1.94 0.365 1.54 0.365 1.54 0.725 1.465 0.725 1.465 0.54 1.46 0.54 1.46 0.41 1.48 0.41 1.48 0.305 2 0.305 2 0.495 2.355 0.495 2.355 0.305 3.36 0.305 3.36 0.79 3.68 0.79 3.68 0.73 3.74 0.73 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 0.895 0.235 0.895 0.235 0.765 0.19 0.765 0.19 0.685 0.56 0.685 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.325 0.885 5.06 0.885 5.06 0.57 5.14 0.57 5.14 0.625 5.325 0.625 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.00305 LAYER Metal1 ;
    ANTENNADIFFAREA 3.7367 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.341775 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.78662875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 67.254773 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.19 1.005 0.72 1.005 0.72 1.055 0.6 1.055 0.6 0.995 0.66 0.995 0.66 0.49 0.72 0.49 0.72 0.79 0.74 0.79 0.74 0.945 1.095 0.945 1.095 0.49 1.19 0.49 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 0 1.77 0 1.65 0.365 1.65 0.365 1.315 0.485 1.315 0.485 1.375 0.425 1.375 0.425 1.65 0.835 1.65 0.835 1.315 0.955 1.315 0.955 1.375 0.895 1.375 0.895 1.65 1.375 1.65 1.375 1.51 1.435 1.51 1.435 1.65 1.775 1.65 1.775 1.51 1.835 1.51 1.835 1.65 2.29 1.65 2.29 1.295 2.35 1.295 2.35 1.65 3.45 1.65 3.45 1.54 3.57 1.54 3.57 1.65 4.165 1.65 4.165 1.54 4.285 1.54 4.285 1.65 5.135 1.65 5.135 1.145 5.195 1.145 5.195 1.65 5.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5.195 0.06 5.195 0.47 5.135 0.47 5.135 0.06 3.52 0.06 3.52 0.47 3.46 0.47 3.46 0.06 2.16 0.06 2.16 0.335 2.22 0.335 2.22 0.395 2.1 0.395 2.1 0.06 1.36 0.06 1.36 0.47 1.3 0.47 1.3 0.06 0.925 0.06 0.925 0.47 0.865 0.47 0.865 0.06 0.51 0.06 0.51 0.585 0.45 0.585 0.45 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.485 1.17 5.34 1.17 5.34 1.045 4.96 1.045 4.96 1.27 4.58 1.27 4.58 1.235 3.84 1.235 3.84 1.195 2.98 1.195 2.98 0.875 2.675 0.875 2.675 0.815 2.98 0.815 2.98 0.65 3.04 0.65 3.04 1.135 3.9 1.135 3.9 1.175 4.58 1.175 4.58 0.855 4.49 0.855 4.49 0.815 4.43 0.815 4.43 0.755 4.55 0.755 4.55 0.795 4.64 0.795 4.64 1.21 4.9 1.21 4.9 0.77 4.96 0.77 4.96 0.985 5.425 0.985 5.425 0.375 5.485 0.375 ;
      POLYGON 4.8 1.11 4.74 1.11 4.74 0.63 3.58 0.63 3.58 0.685 3.46 0.685 3.46 0.57 4.535 0.57 4.535 0.435 4.595 0.435 4.595 0.57 4.8 0.57 ;
      POLYGON 4.48 1.075 4 1.075 4 0.995 4.4 0.995 4.4 0.955 4.48 0.955 ;
      POLYGON 4.48 1.44 3.68 1.44 3.68 1.385 2.61 1.385 2.61 1.195 2.19 1.195 2.19 1.355 1.055 1.355 1.055 1.215 0.25 1.215 0.25 1.31 0.03 1.31 0.03 0.52 0.335 0.52 0.335 0.58 0.09 0.58 0.09 1.155 1.115 1.155 1.115 1.295 2.13 1.295 2.13 1.135 2.67 1.135 2.67 1.325 3.74 1.325 3.74 1.38 4.48 1.38 ;
      POLYGON 4.23 0.895 3.9 0.895 3.9 1.01 3.26 1.01 3.26 1.035 3.14 1.035 3.14 0.525 3.08 0.525 3.08 0.465 3.2 0.465 3.2 0.95 3.84 0.95 3.84 0.835 4.17 0.835 4.17 0.775 4.23 0.775 ;
      POLYGON 2.94 0.525 2.575 0.525 2.575 0.975 2.83 0.975 2.83 1.225 2.77 1.225 2.77 1.035 2.515 1.035 2.515 0.715 2.255 0.715 2.255 0.875 1.8 0.875 1.8 0.73 1.86 0.73 1.86 0.815 2.195 0.815 2.195 0.655 2.515 0.655 2.515 0.465 2.94 0.465 ;
      POLYGON 2.415 1.035 2.03 1.035 2.03 1.195 1.91 1.195 1.91 1.135 1.97 1.135 1.97 1.035 1.6 1.035 1.6 1.095 1.48 1.095 1.48 1.035 1.29 1.035 1.29 0.755 1.35 0.755 1.35 0.975 1.64 0.975 1.64 0.465 1.825 0.465 1.825 0.525 1.7 0.525 1.7 0.975 2.355 0.975 2.355 0.915 2.415 0.915 ;
  END
END DFFRHQX4

MACRO DFFRHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRHQX8 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.54 1.085 6.46 1.085 6.46 1.005 6.465 1.005 6.465 0.605 6.54 0.605 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1074 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.110925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 0.96822175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.44219075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.445 0.81 2.385 0.81 2.385 0.405 1.805 0.405 1.805 0.795 1.66 0.795 1.66 0.6 1.745 0.6 1.745 0.345 2.445 0.345 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.175 0.615 5.965 0.615 5.965 0.705 5.83 0.705 5.83 0.47 6.175 0.47 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.70615 LAYER Metal1 ;
    ANTENNADIFFAREA 4.6892 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.499275 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.4230635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 57.95403325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.63 1.315 0.63 1.315 0.9 1.36 0.9 1.36 1.345 1.3 1.345 1.3 0.96 1.255 0.96 1.255 0.8 0.95 0.8 0.95 1.345 0.89 1.345 0.89 0.73 0.54 0.73 0.54 1.345 0.48 1.345 0.48 0.73 0.13 0.73 0.13 1.345 0.06 1.345 0.06 0.54 0.14 0.54 0.14 0.67 0.49 0.67 0.49 0.54 0.55 0.54 0.55 0.67 0.9 0.67 0.9 0.54 0.96 0.54 0.96 0.74 1.255 0.74 1.255 0.57 1.4 0.57 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 1.77 0 1.77 0 1.65 0.275 1.65 0.275 0.9 0.335 0.9 0.335 1.65 0.685 1.65 0.685 0.9 0.745 0.9 0.745 1.65 1.095 1.65 1.095 0.9 1.155 0.9 1.155 1.65 1.51 1.65 1.51 1.055 1.57 1.055 1.57 1.65 1.955 1.65 1.955 1.25 2.075 1.25 2.075 1.31 2.015 1.31 2.015 1.65 2.46 1.65 2.46 1.25 2.58 1.25 2.58 1.31 2.52 1.31 2.52 1.65 2.955 1.65 2.955 1.54 3.075 1.54 3.075 1.65 3.535 1.65 3.535 1.54 3.655 1.54 3.655 1.65 4.665 1.65 4.665 1.31 4.605 1.31 4.605 1.25 4.725 1.25 4.725 1.65 5.19 1.65 5.19 1.54 5.31 1.54 5.31 1.65 5.95 1.65 5.95 1.185 6.01 1.185 6.01 1.65 6.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 0.06 6.26 0.06 6.26 0.37 6.2 0.37 6.2 0.06 5.955 0.06 5.955 0.31 6.015 0.31 6.015 0.37 5.895 0.37 5.895 0.06 4.87 0.06 4.87 0.32 4.75 0.32 4.75 0.26 4.81 0.26 4.81 0.06 3.46 0.06 3.46 0.17 3.34 0.17 3.34 0.06 2.605 0.06 2.605 0.485 2.545 0.485 2.545 0.06 1.645 0.06 1.645 0.485 1.585 0.485 1.585 0.06 1.165 0.06 1.165 0.485 1.105 0.485 1.105 0.06 0.755 0.06 0.755 0.485 0.695 0.485 0.695 0.06 0.345 0.06 0.345 0.485 0.285 0.485 0.285 0.06 0 0.06 0 -0.06 6.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.53 0.53 6.335 0.53 6.335 1.305 6.275 1.305 6.275 0.865 5.54 0.865 5.54 0.845 5.48 0.845 5.48 0.785 5.6 0.785 5.6 0.805 6.275 0.805 6.275 0.47 6.47 0.47 6.47 0.275 6.53 0.275 ;
      POLYGON 5.73 0.705 5.67 0.705 5.67 0.295 5.22 0.295 5.22 0.715 5.16 0.715 5.16 0.48 4.59 0.48 4.59 0.295 4.27 0.295 4.27 0.67 4.15 0.67 4.15 0.61 4.21 0.61 4.21 0.295 3.89 0.295 3.89 0.99 3.1 0.99 3.1 0.63 3.04 0.63 3.04 0.57 3.16 0.57 3.16 0.93 3.83 0.93 3.83 0.235 4.65 0.235 4.65 0.42 5.16 0.42 5.16 0.235 5.73 0.235 ;
      POLYGON 5.7 1.23 5.64 1.23 5.64 1.025 5.32 1.025 5.32 0.935 4.585 0.935 4.585 0.74 4.645 0.74 4.645 0.875 5.32 0.875 5.32 0.395 5.44 0.395 5.44 0.455 5.38 0.455 5.38 0.965 5.7 0.965 ;
      POLYGON 5.59 1.39 5.47 1.39 5.47 1.365 4.825 1.365 4.825 1.15 4.205 1.15 4.205 0.77 4.325 0.77 4.325 0.83 4.265 0.83 4.265 1.09 4.885 1.09 4.885 1.305 5.53 1.305 5.53 1.33 5.59 1.33 ;
      POLYGON 5.525 1.205 4.985 1.205 4.985 1.085 5.065 1.085 5.065 1.125 5.525 1.125 ;
      POLYGON 5.04 0.775 4.98 0.775 4.98 0.64 4.485 0.64 4.485 0.99 4.365 0.99 4.365 0.93 4.425 0.93 4.425 0.64 4.37 0.64 4.37 0.395 4.49 0.395 4.49 0.58 5.04 0.58 ;
      RECT 2.66 1.38 4.45 1.44 ;
      POLYGON 4.11 0.455 4.05 0.455 4.05 1.15 2.065 1.15 2.065 0.74 2.125 0.74 2.125 1.09 2.94 1.09 2.94 0.85 2.91 0.85 2.91 0.73 3 0.73 3 1.09 3.99 1.09 3.99 0.395 4.11 0.395 ;
      POLYGON 3.73 0.815 3.26 0.815 3.26 0.735 3.65 0.735 3.65 0.55 3.73 0.55 ;
      POLYGON 3.55 0.625 3.26 0.625 3.26 0.47 2.915 0.47 2.915 0.63 2.81 0.63 2.81 0.93 2.84 0.93 2.84 0.99 2.225 0.99 2.225 0.64 1.965 0.64 1.965 0.955 1.84 0.955 1.84 1.34 1.78 1.34 1.78 0.955 1.475 0.955 1.475 0.805 1.415 0.805 1.415 0.745 1.535 0.745 1.535 0.895 1.905 0.895 1.905 0.58 1.985 0.58 1.985 0.505 2.045 0.505 2.045 0.58 2.285 0.58 2.285 0.93 2.75 0.93 2.75 0.57 2.855 0.57 2.855 0.41 3.32 0.41 3.32 0.565 3.55 0.565 ;
  END
END DFFRHQX8

MACRO DFFRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRX1 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.32595 LAYER Metal1 ;
    ANTENNADIFFAREA 2.408925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2205 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.548526 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 84.2312925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.73 0.585 0.69 0.585 0.69 1.455 0.63 1.455 0.63 0.73 0.61 0.73 0.61 0.6 0.63 0.6 0.63 0.515 0.67 0.515 0.67 0.325 0.73 0.325 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.32595 LAYER Metal1 ;
    ANTENNADIFFAREA 2.408925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2205 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.548526 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 84.2312925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.05 0.4 0.13 1.29 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0687 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.12037025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 25.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.355 0.775 1.605 0.895 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.24074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.79 0.855 1.03 1.06 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.43 0.635 3.555 0.87 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 0 1.77 0 1.65 0.305 1.65 0.305 1.285 0.365 1.285 0.365 1.65 0.865 1.65 0.865 1.51 0.925 1.51 0.925 1.65 1.285 1.65 1.285 1.505 1.345 1.505 1.345 1.65 1.655 1.65 1.655 1.54 1.775 1.54 1.775 1.65 2.36 1.65 2.36 1.54 2.48 1.54 2.48 1.65 2.79 1.65 2.79 1.51 2.85 1.51 2.85 1.65 3.5 1.65 3.5 1.51 3.56 1.51 3.56 1.65 4 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.46 0.06 3.46 0.555 3.4 0.555 3.4 0.06 2.525 0.06 2.525 0.45 2.465 0.45 2.465 0.06 1.715 0.06 1.715 0.475 1.655 0.475 1.655 0.06 0.935 0.06 0.935 0.56 0.875 0.56 0.875 0.06 0.365 0.06 0.365 0.335 0.305 0.335 0.305 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.795 1.195 3.735 1.195 3.735 1 3.34 1 3.34 1.035 3.28 1.035 3.28 0.36 2.74 0.36 2.74 0.59 2.345 0.59 2.345 0.3 2.155 0.3 2.155 0.675 2.005 0.675 2.005 0.885 1.945 0.885 1.945 0.615 2.095 0.615 2.095 0.185 2.155 0.185 2.155 0.24 2.405 0.24 2.405 0.53 2.675 0.53 2.675 0.3 3.34 0.3 3.34 0.94 3.62 0.94 3.62 0.46 3.68 0.46 3.68 0.94 3.795 0.94 ;
      POLYGON 3.76 1.42 2.81 1.42 2.81 1.28 1.03 1.28 1.03 1.16 1.115 1.16 1.115 0.465 1.175 0.465 1.175 1.22 2.105 1.22 2.105 0.765 2.165 0.765 2.165 1.22 2.87 1.22 2.87 1.36 3.76 1.36 ;
      POLYGON 3.275 1.255 3.215 1.255 3.215 1.195 3.15 1.195 3.15 0.87 2.425 0.87 2.425 0.895 2.365 0.895 2.365 0.775 2.425 0.775 2.425 0.81 3.01 0.81 3.01 0.46 3.07 0.46 3.07 0.81 3.21 0.81 3.21 1.135 3.275 1.135 ;
      POLYGON 3.07 1.195 3.01 1.195 3.01 1.1 2.595 1.1 2.595 1.04 3.07 1.04 ;
      POLYGON 2.855 0.71 2.285 0.71 2.285 1.09 2.225 1.09 2.225 0.38 2.285 0.38 2.285 0.65 2.855 0.65 ;
      RECT 1.495 1.38 2.64 1.44 ;
      POLYGON 2.035 0.5 1.885 0.5 1.885 0.965 2.035 0.965 2.035 1.115 1.975 1.115 1.975 1.025 1.825 1.025 1.825 0.685 1.385 0.685 1.385 0.565 1.445 0.565 1.445 0.625 1.825 0.625 1.825 0.44 1.975 0.44 1.975 0.375 2.035 0.375 ;
      POLYGON 1.765 1.12 1.235 1.12 1.235 0.385 1.055 0.385 1.055 0.715 0.77 0.715 0.77 0.655 0.995 0.655 0.995 0.32 1.295 0.32 1.295 0.385 1.44 0.385 1.44 0.445 1.295 0.445 1.295 1.06 1.705 1.06 1.705 0.775 1.765 0.775 ;
      POLYGON 0.53 1.02 0.47 1.02 0.47 0.83 0.19 0.83 0.19 0.77 0.47 0.77 0.47 0.54 0.53 0.54 ;
  END
END DFFRX1

MACRO DFFRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRX2 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.588 LAYER Metal1 ;
    ANTENNADIFFAREA 2.74135 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.285975 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.049742 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 72.1321795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.965 1.11 3.895 1.11 3.895 1.305 3.835 1.305 3.835 0.975 3.785 0.975 3.785 0.565 3.925 0.565 3.925 0.625 3.845 0.625 3.845 0.915 3.965 0.915 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.588 LAYER Metal1 ;
    ANTENNADIFFAREA 2.74135 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.285975 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.049742 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 72.1321795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.5 1.11 3.48 1.11 3.48 1.305 3.42 1.305 3.42 0.535 3.48 0.535 3.48 0.925 3.5 0.925 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.425926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.32 1.085 3.06 1.085 3.06 0.89 3.12 0.89 3.12 1.005 3.32 1.005 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.039375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.80952375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.605 0.935 1.225 0.935 1.225 0.815 1.355 0.815 1.355 0.855 1.605 0.855 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.445 1.185 0.235 1.185 0.235 1.005 0.365 1.005 0.365 0.815 0.445 0.815 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.34 1.65 0.34 1.51 0.4 1.51 0.4 1.65 0.965 1.65 0.965 1.54 1.085 1.54 1.085 1.65 1.465 1.65 1.465 1.43 1.525 1.43 1.525 1.65 2.405 1.65 2.405 1.51 2.465 1.51 2.465 1.65 2.83 1.65 2.83 1.51 2.89 1.51 2.89 1.65 3.175 1.65 3.175 1.185 3.235 1.185 3.235 1.65 3.625 1.65 3.625 0.925 3.685 0.925 3.685 1.65 4.04 1.65 4.04 1.01 4.1 1.01 4.1 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 4.16 0.06 4.16 0.17 4.04 0.17 4.04 0.06 3.745 0.06 3.745 0.17 3.625 0.17 3.625 0.06 3.24 0.06 3.24 0.63 3.18 0.63 3.18 0.06 2.435 0.06 2.435 0.585 2.375 0.585 2.375 0.06 1.505 0.06 1.505 0.425 1.445 0.425 1.445 0.06 0.57 0.06 0.57 0.495 0.63 0.495 0.63 0.555 0.51 0.555 0.51 0.06 0.37 0.06 0.37 0.555 0.31 0.555 0.31 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.305 1.035 4.245 1.035 4.245 0.785 3.945 0.785 3.945 0.725 4.245 0.725 4.245 0.535 4.305 0.535 ;
      POLYGON 4.26 0.43 3.825 0.43 3.825 0.435 3.61 0.435 3.61 0.825 3.55 0.825 3.55 0.435 3.36 0.435 3.36 0.85 3.26 0.85 3.26 0.79 3.06 0.79 3.06 0.425 2.76 0.425 2.76 0.525 2.865 0.525 2.865 0.88 2.655 0.88 2.655 1.095 2.595 1.095 2.595 0.88 2.41 0.88 2.41 0.935 2.35 0.935 2.35 0.815 2.805 0.815 2.805 0.585 2.7 0.585 2.7 0.365 3.12 0.365 3.12 0.73 3.3 0.73 3.3 0.375 3.79 0.375 3.79 0.37 4.26 0.37 ;
      POLYGON 3.03 1.35 0.14 1.35 0.14 1.29 2.94 1.29 2.94 0.535 3 0.535 3 1.185 3.03 1.185 ;
      POLYGON 2.725 0.745 2.29 0.745 2.29 1.125 2.035 1.125 2.035 1.065 2.23 1.065 2.23 0.745 1.965 0.745 1.965 0.49 2.025 0.49 2.025 0.685 2.725 0.685 ;
      POLYGON 2.17 0.955 2.11 0.955 2.11 0.89 1.83 0.89 1.83 0.39 1.635 0.39 1.635 0.565 1.255 0.565 1.255 0.395 0.79 0.395 0.79 0.715 0.605 0.715 0.605 0.9 0.545 0.9 0.545 0.715 0.165 0.715 0.165 1.095 0.105 1.095 0.105 0.46 0.165 0.46 0.165 0.655 0.73 0.655 0.73 0.335 0.955 0.335 0.955 0.265 1.075 0.265 1.075 0.335 1.315 0.335 1.315 0.505 1.575 0.505 1.575 0.33 1.89 0.33 1.89 0.83 2.17 0.83 ;
      POLYGON 1.76 1.19 1.7 1.19 1.7 1.055 1.075 1.055 1.075 0.9 1.135 0.9 1.135 0.995 1.7 0.995 1.7 0.49 1.76 0.49 ;
      POLYGON 1.62 0.77 1.56 0.77 1.56 0.71 0.95 0.71 0.95 0.97 0.765 0.97 0.765 1.09 0.63 1.09 0.63 1.03 0.705 1.03 0.705 0.91 0.89 0.91 0.89 0.495 1.01 0.495 1.01 0.555 0.95 0.555 0.95 0.65 1.62 0.65 ;
      POLYGON 1.32 1.19 0.865 1.19 0.865 1.07 0.925 1.07 0.925 1.12 1.32 1.12 ;
  END
END DFFRX2

MACRO DFFRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRX4 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.21365 LAYER Metal1 ;
    ANTENNADIFFAREA 3.69945 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4392 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.31705375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 56.420765 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.06 0.63 4.605 0.63 4.605 1.05 4.99 1.05 4.99 1.33 4.93 1.33 4.93 1.11 4.58 1.11 4.58 1.33 4.52 1.33 4.52 1.11 4.435 1.11 4.435 0.98 4.53 0.98 4.53 0.57 5.06 0.57 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.21365 LAYER Metal1 ;
    ANTENNADIFFAREA 3.69945 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4392 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.31705375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 56.420765 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.18 0.61 3.785 0.61 3.785 0.79 3.965 0.79 3.965 0.94 4.15 0.94 4.15 1.33 4.09 1.33 4.09 1 3.74 1 3.74 1.33 3.68 1.33 3.68 0.94 3.725 0.94 3.725 0.61 3.59 0.61 3.59 0.55 4.18 0.55 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06255 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 12.82973625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.37 0.63 2.775 0.63 2.775 0.47 2.485 0.47 2.485 0.38 1.96 0.38 1.96 0.91 1.575 0.91 1.575 0.85 1.9 0.85 1.9 0.735 1.86 0.735 1.86 0.6 1.9 0.6 1.9 0.32 2.545 0.32 2.545 0.41 2.835 0.41 2.835 0.57 3.37 0.57 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.462963 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.81 0.865 0.74 0.865 0.74 1.2 0.66 1.2 0.66 0.785 0.81 0.785 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.9814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.205 0.92 0.035 0.92 0.035 0.79 0.125 0.79 0.125 0.605 0.205 0.605 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.12 0.13 1.12 0.13 1.65 0.665 1.65 0.665 1.51 0.725 1.51 0.725 1.65 1.3 1.65 1.3 1.54 1.42 1.54 1.42 1.65 1.795 1.65 1.795 1.54 1.915 1.54 1.915 1.65 2.57 1.65 2.57 1.115 2.63 1.115 2.63 1.65 3.045 1.65 3.045 1.085 3.105 1.085 3.105 1.65 3.455 1.65 3.455 1.21 3.515 1.21 3.515 1.65 3.885 1.65 3.885 1.1 3.945 1.1 3.945 1.65 4.295 1.65 4.295 0.94 4.355 0.94 4.355 1.65 4.725 1.65 4.725 1.21 4.785 1.21 4.785 1.65 5.135 1.65 5.135 1.08 5.195 1.08 5.195 1.65 5.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5.3 0.06 5.3 0.52 5.24 0.52 5.24 0.06 4.885 0.06 4.885 0.17 4.765 0.17 4.765 0.06 4.415 0.06 4.415 0.17 4.295 0.17 4.295 0.06 3.945 0.06 3.945 0.17 3.825 0.17 3.825 0.06 3.475 0.06 3.475 0.17 3.355 0.17 3.355 0.06 2.765 0.06 2.765 0.17 2.645 0.17 2.645 0.06 1.81 0.06 1.81 0.43 1.78 0.43 1.78 0.555 1.72 0.555 1.72 0.06 0.93 0.06 0.93 0.465 0.99 0.465 0.99 0.525 0.87 0.525 0.87 0.06 0.71 0.06 0.71 0.465 0.77 0.465 0.77 0.525 0.65 0.525 0.65 0.06 0.17 0.06 0.17 0.265 0.11 0.265 0.11 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.505 0.68 5.455 0.68 5.455 0.98 5.4 0.98 5.4 1.33 5.34 1.33 5.34 0.98 5.055 0.98 5.055 0.8 5.175 0.8 5.175 0.92 5.395 0.92 5.395 0.62 5.445 0.62 5.445 0.54 5.505 0.54 ;
      POLYGON 5.335 0.82 5.275 0.82 5.275 0.7 5.12 0.7 5.12 0.44 4.34 0.44 4.34 0.77 4.28 0.77 4.28 0.83 4.22 0.83 4.22 0.71 4.28 0.71 4.28 0.44 3.015 0.44 3.015 0.38 5.18 0.38 5.18 0.64 5.335 0.64 ;
      POLYGON 3.58 0.95 3.31 0.95 3.31 1.33 3.25 1.33 3.25 0.95 2.9 0.95 2.9 1.33 2.84 1.33 2.84 0.95 2.475 0.95 2.475 0.89 3.52 0.89 3.52 0.78 3.58 0.78 ;
      POLYGON 3.005 0.79 2.535 0.79 2.535 0.63 2.27 0.63 2.27 1.14 2.21 1.14 2.21 0.57 2.225 0.57 2.225 0.46 2.285 0.46 2.285 0.57 2.595 0.57 2.595 0.73 3.005 0.73 ;
      POLYGON 2.415 1.37 0.6 1.37 0.6 1.43 0.54 1.43 0.54 1.37 0.275 1.37 0.275 0.46 0.335 0.46 0.335 1.31 2.355 1.31 2.355 0.7 2.415 0.7 ;
      POLYGON 2.08 1.03 2.065 1.03 2.065 1.165 2.005 1.165 2.005 1.03 1.42 1.03 1.42 0.85 1.48 0.85 1.48 0.97 2.02 0.97 2.02 0.46 2.08 0.46 ;
      POLYGON 1.78 0.775 1.72 0.775 1.72 0.675 1.27 0.675 1.27 0.985 1.15 0.985 1.15 1.11 1.065 1.11 1.065 1.17 1.005 1.17 1.005 1.05 1.09 1.05 1.09 0.925 1.21 0.925 1.21 0.49 1.33 0.49 1.33 0.55 1.27 0.55 1.27 0.615 1.78 0.615 ;
      POLYGON 1.68 1.21 1.21 1.21 1.21 1.085 1.27 1.085 1.27 1.12 1.68 1.12 ;
      POLYGON 1.63 0.28 1.115 0.28 1.115 0.685 0.97 0.685 0.97 0.89 1.03 0.89 1.03 0.95 0.91 0.95 0.91 0.685 0.535 0.685 0.535 1.145 0.475 1.145 0.475 0.46 0.535 0.46 0.535 0.625 1.055 0.625 1.055 0.22 1.57 0.22 1.57 0.145 1.63 0.145 ;
  END
END DFFRX4

MACRO DFFRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRXL 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.67995 LAYER Metal1 ;
    ANTENNADIFFAREA 2.792975 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1944 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.785751 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 105.67901225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.555 0.885 0.555 0.885 0.98 0.94 0.98 0.94 1.11 0.885 1.11 0.885 1.22 0.825 1.22 0.825 0.495 0.94 0.495 0.94 0.435 1 0.435 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.67995 LAYER Metal1 ;
    ANTENNADIFFAREA 2.792975 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1944 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.785751 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 105.67901225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.29 1.02 0.21 1.02 0.21 0.73 0.06 0.73 0.06 0.6 0.21 0.6 0.21 0.54 0.29 0.54 ;
    END
  END QN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.09 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.77777775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 34.25925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.785 0.72 2.125 0.96 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 0.895 1.315 0.895 1.315 1.265 1.235 1.265 1.235 0.815 1.365 0.815 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.435 0.625 4.655 0.815 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 1.77 0 1.77 0 1.65 0.49 1.65 0.49 1.285 0.55 1.285 0.55 1.65 1.06 1.65 1.06 1.51 1.12 1.51 1.12 1.65 1.805 1.65 1.805 1.51 1.865 1.51 1.865 1.65 2.175 1.65 2.175 1.54 2.295 1.54 2.295 1.65 3.235 1.65 3.235 1.54 3.355 1.54 3.355 1.65 3.615 1.65 3.615 1.51 3.675 1.51 3.675 1.65 4.635 1.65 4.635 1.51 4.695 1.51 4.695 1.65 5 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 0.06 4.555 0.06 4.555 0.525 4.435 0.525 4.435 0.465 4.495 0.465 4.495 0.06 3.5 0.06 3.5 0.25 3.38 0.25 3.38 0.19 3.44 0.19 3.44 0.06 2.235 0.06 2.235 0.455 2.175 0.455 2.175 0.06 1.205 0.06 1.205 0.55 1.145 0.55 1.145 0.06 0.52 0.06 0.52 0.635 0.46 0.635 0.46 0.06 0 0.06 0 -0.06 5 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.96 1 4.755 1 4.755 0.975 4.335 0.975 4.335 1.035 4.275 1.035 4.275 0.36 3.66 0.36 3.66 0.41 3.22 0.41 3.22 0.385 2.9 0.385 2.9 0.715 2.605 0.715 2.605 0.875 2.545 0.875 2.545 0.655 2.84 0.655 2.84 0.325 3.28 0.325 3.28 0.35 3.6 0.35 3.6 0.3 4.335 0.3 4.335 0.915 4.755 0.915 4.755 0.46 4.815 0.46 4.815 0.94 4.96 0.94 ;
      POLYGON 4.865 1.285 4.805 1.285 4.805 1.225 4.535 1.225 4.535 1.415 4.11 1.415 4.11 1.42 3.99 1.42 3.99 1.415 3.775 1.415 3.775 1.41 3.615 1.41 3.615 1.28 1.415 1.28 1.415 1.1 1.465 1.1 1.465 0.54 1.525 0.54 1.525 1.22 2.78 1.22 2.78 0.875 2.82 0.875 2.82 0.815 2.88 0.815 2.88 0.935 2.84 0.935 2.84 1.22 3.675 1.22 3.675 1.35 3.835 1.35 3.835 1.355 4.475 1.355 4.475 1.165 4.865 1.165 ;
      POLYGON 4.22 1.255 4.16 1.255 4.16 1.195 4.115 1.195 4.115 0.87 3.16 0.87 3.16 0.81 3.93 0.81 3.93 0.46 3.99 0.46 3.99 0.81 4.175 0.81 4.175 1.135 4.22 1.135 ;
      POLYGON 4.015 1.195 3.935 1.195 3.935 1.12 3.515 1.12 3.515 1.04 4.015 1.04 ;
      POLYGON 3.775 0.71 3.06 0.71 3.06 1.095 2.94 1.095 2.94 1.035 3 1.035 3 0.485 3.12 0.485 3.12 0.65 3.775 0.65 ;
      RECT 2.015 1.38 3.515 1.44 ;
      POLYGON 2.74 0.545 2.445 0.545 2.445 1.005 2.665 1.005 2.665 1.065 2.385 1.065 2.385 0.62 1.865 0.62 1.865 0.56 2.385 0.56 2.385 0.485 2.74 0.485 ;
      POLYGON 2.285 1.12 1.625 1.12 1.625 0.4 1.82 0.4 1.82 0.3 1.365 0.3 1.365 0.715 0.985 0.715 0.985 0.655 1.305 0.655 1.305 0.24 1.88 0.24 1.88 0.46 1.685 0.46 1.685 1.06 2.225 1.06 2.225 0.815 2.285 0.815 ;
      POLYGON 0.725 1.02 0.645 1.02 0.645 0.815 0.39 0.815 0.39 0.735 0.645 0.735 0.645 0.54 0.725 0.54 ;
  END
END DFFRXL

MACRO DFFSHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSHQX1 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.186775 LAYER Metal1 ;
    ANTENNADIFFAREA 2.329325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.23085 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.4727095 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 75.77647825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.14 0.74 0.13 0.74 0.13 1.29 0.07 1.29 0.07 0.74 0.06 0.74 0.06 0.6 0.07 0.6 0.07 0.54 0.13 0.54 0.13 0.6 0.14 0.6 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.29629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.545 0.775 3.74 0.92 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.184466 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.565 1.11 3.335 1.11 3.335 0.785 3.415 0.785 3.415 0.98 3.565 0.98 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 16.21359225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.25 0.82 2.19 0.82 2.19 0.75 2.02 0.75 2.02 0.41 1.11 0.41 1.11 0.97 0.795 0.97 0.795 0.91 1.05 0.91 1.05 0.625 1.03 0.625 1.03 0.545 1.05 0.545 1.05 0.35 2.08 0.35 2.08 0.69 2.25 0.69 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 1.77 0 1.77 0 1.65 0.275 1.65 0.275 0.93 0.335 0.93 0.335 1.65 0.685 1.65 0.685 1.36 0.745 1.36 0.745 1.65 1.065 1.65 1.065 1.39 1.185 1.39 1.185 1.45 1.125 1.45 1.125 1.65 2.17 1.65 2.17 1.54 2.29 1.54 2.29 1.65 2.695 1.65 2.695 1.215 2.755 1.215 2.755 1.65 3.41 1.65 3.41 1.345 3.47 1.345 3.47 1.65 3.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 0.06 3.525 0.06 3.525 0.535 3.465 0.535 3.465 0.06 2.755 0.06 2.755 0.385 2.815 0.385 2.815 0.445 2.695 0.445 2.695 0.06 2.2 0.06 2.2 0.61 2.14 0.61 2.14 0.06 0.745 0.06 0.745 0.565 0.685 0.565 0.685 0.06 0.335 0.06 0.335 0.52 0.275 0.52 0.275 0.06 0 0.06 0 -0.06 3.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.73 0.695 3.28 0.695 3.28 0.725 3.26 0.725 3.26 1.225 3.71 1.225 3.71 1.37 3.65 1.37 3.65 1.285 3.26 1.285 3.26 1.435 3.02 1.435 3.02 1.475 2.9 1.475 2.9 1.115 2.635 1.115 2.635 1.44 2.01 1.44 2.01 1.38 2.575 1.38 2.575 1.055 2.96 1.055 2.96 1.375 3.2 1.375 3.2 0.635 3.22 0.635 3.22 0.585 3.28 0.585 3.28 0.635 3.67 0.635 3.67 0.44 3.73 0.44 ;
      POLYGON 3.14 1.275 3.08 1.275 3.08 0.925 2.575 0.925 2.575 0.865 3.08 0.865 3.08 0.44 3.14 0.44 ;
      POLYGON 3.02 0.73 2.96 0.73 2.96 0.605 2.57 0.605 2.57 0.435 2.39 0.435 2.39 0.96 1.995 0.96 1.995 1.06 2.055 1.06 2.055 1.12 1.935 1.12 1.935 0.96 1.9 0.96 1.9 0.49 1.96 0.49 1.96 0.9 2.33 0.9 2.33 0.375 2.63 0.375 2.63 0.545 3.02 0.545 ;
      POLYGON 2.86 0.765 2.515 0.765 2.515 1.28 1.825 1.28 1.825 1.35 1.765 1.35 1.765 0.74 1.58 0.74 1.58 0.56 1.7 0.56 1.7 0.68 1.825 0.68 1.825 1.22 2.45 1.22 2.45 0.52 2.51 0.52 2.51 0.705 2.86 0.705 ;
      POLYGON 1.68 0.96 1.305 0.96 1.305 0.84 1.385 0.84 1.385 0.88 1.68 0.88 ;
      POLYGON 1.605 1.35 1.545 1.35 1.545 1.13 0.635 1.13 0.635 1.01 0.695 1.01 0.695 1.07 1.17 1.07 1.17 0.56 1.48 0.56 1.48 0.62 1.23 0.62 1.23 1.07 1.605 1.07 ;
      POLYGON 1.4 1.35 1.34 1.35 1.34 1.29 0.95 1.29 0.95 1.35 0.89 1.35 0.89 1.23 1.4 1.23 ;
      POLYGON 0.99 0.81 0.535 0.81 0.535 1.48 0.475 1.48 0.475 0.77 0.29 0.77 0.29 0.83 0.23 0.83 0.23 0.71 0.48 0.71 0.48 0.53 0.54 0.53 0.54 0.75 0.93 0.75 0.93 0.69 0.99 0.69 ;
  END
END DFFSHQX1

MACRO DFFSHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSHQX2 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5684 LAYER Metal1 ;
    ANTENNADIFFAREA 2.83185 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2601 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.8746635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 76.793541 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.54 0.34 1.29 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.77 0.985 4.635 0.985 4.635 0.79 4.465 0.79 4.465 0.71 4.77 0.71 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.0841425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.235 0.71 4.365 1.05 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 17.9288025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.94 0.82 2.88 0.82 2.88 0.705 2.66 0.705 2.66 0.41 1.52 0.41 1.52 0.6 1.54 0.6 1.54 0.73 1.52 0.73 1.52 0.92 1.17 0.92 1.17 0.86 1.46 0.86 1.46 0.35 2.72 0.35 2.72 0.645 2.94 0.645 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.075 1.65 0.075 0.9 0.135 0.9 0.135 1.65 0.485 1.65 0.485 0.93 0.545 0.93 0.545 1.65 1.055 1.65 1.055 1.31 1.115 1.31 1.115 1.65 1.435 1.65 1.435 1.34 1.555 1.34 1.555 1.4 1.495 1.4 1.495 1.65 2.895 1.65 2.895 1.54 3.015 1.54 3.015 1.65 3.52 1.65 3.52 1.15 3.58 1.15 3.58 1.65 4.34 1.65 4.34 1.31 4.4 1.31 4.4 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 4.41 0.06 4.41 0.45 4.35 0.45 4.35 0.06 3.58 0.06 3.58 0.17 3.46 0.17 3.46 0.06 2.88 0.06 2.88 0.485 2.94 0.485 2.94 0.545 2.82 0.545 2.82 0.06 1.115 0.06 1.115 0.515 1.055 0.515 1.055 0.06 0.545 0.06 0.545 0.52 0.485 0.52 0.485 0.06 0.135 0.06 0.135 0.52 0.075 0.52 0.075 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.615 0.61 4.135 0.61 4.135 1.15 4.615 1.15 4.615 1.335 4.555 1.335 4.555 1.21 4.135 1.21 4.135 1.4 3.735 1.4 3.735 1.05 3.42 1.05 3.42 1.37 2.735 1.37 2.735 1.31 3.36 1.31 3.36 0.99 3.795 0.99 3.795 1.34 4.075 1.34 4.075 0.55 4.555 0.55 4.555 0.355 4.615 0.355 ;
      POLYGON 3.975 1.24 3.915 1.24 3.915 0.82 3.36 0.82 3.36 0.76 3.915 0.76 3.915 0.355 3.975 0.355 ;
      POLYGON 3.815 0.645 3.755 0.645 3.755 0.44 3.1 0.44 3.1 1.05 2.5 1.05 2.5 0.79 2.4 0.79 2.4 0.67 2.5 0.67 2.5 0.57 2.44 0.57 2.44 0.51 2.56 0.51 2.56 0.99 3.04 0.99 3.04 0.38 3.815 0.38 ;
      POLYGON 3.655 0.66 3.26 0.66 3.26 1.21 2.3 1.21 2.3 1.3 2.24 1.3 2.24 0.57 2.005 0.57 2.005 0.51 2.3 0.51 2.3 1.15 3.2 1.15 3.2 0.54 3.26 0.54 3.26 0.6 3.655 0.6 ;
      POLYGON 2.14 0.92 2.06 0.92 2.06 0.8 1.8 0.8 1.8 0.68 1.88 0.68 1.88 0.72 2.14 0.72 ;
      POLYGON 2.095 1.3 2.035 1.3 2.035 1.08 1.01 1.08 1.01 0.96 1.07 0.96 1.07 1.02 1.64 1.02 1.64 0.51 1.875 0.51 1.875 0.57 1.7 0.57 1.7 1.02 2.095 1.02 ;
      POLYGON 1.89 1.3 1.83 1.3 1.83 1.24 1.32 1.24 1.32 1.3 1.26 1.3 1.26 1.18 1.89 1.18 ;
      POLYGON 1.36 0.76 0.91 0.76 0.91 1.43 0.85 1.43 0.85 0.77 0.5 0.77 0.5 0.83 0.44 0.83 0.44 0.71 0.85 0.71 0.85 0.48 0.91 0.48 0.91 0.7 1.3 0.7 1.3 0.64 1.36 0.64 ;
  END
END DFFSHQX2

MACRO DFFSHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSHQX4 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.365 0.895 5.235 0.895 5.235 0.815 5.285 0.815 5.285 0.445 5.365 0.445 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.785 0.895 4.385 0.895 4.385 0.715 4.465 0.715 4.465 0.815 4.785 0.815 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 16.21359225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.075 0.7 3.015 0.7 3.015 0.575 2.75 0.575 2.75 0.415 1.92 0.415 1.92 0.6 1.94 0.6 1.94 0.73 1.92 0.73 1.92 0.925 1.445 0.925 1.445 0.865 1.86 0.865 1.86 0.355 2.81 0.355 2.81 0.515 3.075 0.515 ;
    END
  END SN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.094525 LAYER Metal1 ;
    ANTENNADIFFAREA 3.324925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.341775 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.0542755 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 70.520079 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.775 1.465 0.715 1.465 0.715 0.73 0.365 0.73 0.365 1.465 0.305 1.465 0.305 0.73 0.26 0.73 0.26 0.6 0.305 0.6 0.305 0.54 0.365 0.54 0.365 0.67 0.715 0.67 0.715 0.54 0.775 0.54 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 0 1.77 0 1.65 0.1 1.65 0.1 1.075 0.16 1.075 0.16 1.65 0.51 1.65 0.51 1.075 0.57 1.075 0.57 1.65 0.92 1.65 0.92 1.155 0.98 1.155 0.98 1.65 1.35 1.65 1.35 1.185 1.41 1.185 1.41 1.65 1.81 1.65 1.81 1.345 1.87 1.345 1.87 1.65 2.995 1.65 2.995 1.54 3.115 1.54 3.115 1.65 3.465 1.65 3.465 1.54 3.585 1.54 3.585 1.65 4.47 1.65 4.47 1.155 4.53 1.155 4.53 1.65 5.35 1.65 5.35 0.995 5.41 0.995 5.41 1.65 5.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5.525 0.06 5.525 0.635 5.465 0.635 5.465 0.06 4.465 0.06 4.465 0.395 4.525 0.395 4.525 0.455 4.405 0.455 4.405 0.06 3.805 0.06 3.805 0.485 3.745 0.485 3.745 0.06 3.03 0.06 3.03 0.415 2.91 0.415 2.91 0.355 2.97 0.355 2.97 0.06 1.39 0.06 1.39 0.52 1.33 0.52 1.33 0.06 0.98 0.06 0.98 0.52 0.92 0.52 0.92 0.06 0.57 0.06 0.57 0.52 0.51 0.52 0.51 0.06 0.16 0.06 0.16 0.52 0.1 0.52 0.1 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.235 1.055 5.075 1.055 5.075 0.655 5.125 0.655 5.125 0.38 4.685 0.38 4.685 0.715 4.565 0.715 4.565 0.615 4.28 0.615 4.28 0.7 4.125 0.7 4.125 1.215 2.635 1.215 2.635 0.895 2.26 0.895 2.26 0.76 2.2 0.76 2.2 0.7 2.32 0.7 2.32 0.835 2.755 0.835 2.755 0.895 2.695 0.895 2.695 1.155 4.065 1.155 4.065 0.83 3.875 0.83 3.875 0.77 4.065 0.77 4.065 0.555 4.625 0.555 4.625 0.32 5.185 0.32 5.185 0.715 5.135 0.715 5.135 0.995 5.235 0.995 ;
      POLYGON 5.005 0.54 4.945 0.54 4.945 1.18 4.725 1.18 4.725 1.055 4.285 1.055 4.285 1.415 2.37 1.415 2.37 1.355 4.225 1.355 4.225 0.805 4.285 0.805 4.285 0.995 4.885 0.995 4.885 0.48 5.005 0.48 ;
      POLYGON 4.215 0.455 3.965 0.455 3.965 0.645 3.775 0.645 3.775 0.995 3.965 0.995 3.965 1.055 3.715 1.055 3.715 0.86 3.335 0.86 3.335 0.73 3.395 0.73 3.395 0.8 3.715 0.8 3.715 0.585 3.905 0.585 3.905 0.395 4.215 0.395 ;
      POLYGON 3.615 0.7 3.495 0.7 3.495 0.63 3.235 0.63 3.235 0.96 3.35 0.96 3.35 1.02 3.175 1.02 3.175 0.86 2.915 0.86 2.915 1.055 2.795 1.055 2.795 0.995 2.855 0.995 2.855 0.735 2.505 0.735 2.505 0.575 2.445 0.575 2.445 0.515 2.565 0.515 2.565 0.675 2.915 0.675 2.915 0.8 3.175 0.8 3.175 0.57 3.25 0.57 3.25 0.41 3.31 0.41 3.31 0.57 3.555 0.57 3.555 0.64 3.615 0.64 ;
      POLYGON 2.535 1.255 2.475 1.255 2.475 1.085 1.285 1.085 1.285 0.965 1.345 0.965 1.345 1.025 2.04 1.025 2.04 0.515 2.29 0.515 2.29 0.575 2.1 0.575 2.1 1.025 2.535 1.025 ;
      POLYGON 2.36 1.245 1.665 1.245 1.665 1.465 1.605 1.465 1.605 1.185 2.36 1.185 ;
      POLYGON 1.73 0.765 1.185 0.765 1.185 1.465 1.125 1.465 1.125 0.76 0.935 0.76 0.935 0.82 0.875 0.82 0.875 0.7 1.125 0.7 1.125 0.485 1.185 0.485 1.185 0.705 1.67 0.705 1.67 0.645 1.73 0.645 ;
  END
END DFFSHQX4

MACRO DFFSHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSHQX8 0 0 ;
  SIZE 6.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.17 0.98 5.87 0.98 5.87 0.9 6.035 0.9 6.035 0.7 6.17 0.7 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.77 0.98 5.47 0.98 5.47 0.815 5.69 0.815 5.69 0.7 5.77 0.7 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 16.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.085 0.73 4.025 0.73 4.025 0.33 3.805 0.33 3.805 0.295 2.92 0.295 2.92 0.41 2.94 0.41 2.94 0.54 2.92 0.54 2.92 0.855 2.585 0.855 2.585 0.795 2.86 0.795 2.86 0.235 3.865 0.235 3.865 0.27 4.085 0.27 ;
    END
  END SN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.313575 LAYER Metal1 ;
    ANTENNADIFFAREA 4.00885 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.499275 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.63677325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 51.59080675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.37 1.345 1.31 1.345 1.31 0.66 0.96 0.66 0.96 1.345 0.9 1.345 0.9 0.66 0.55 0.66 0.55 1.345 0.49 1.345 0.49 0.66 0.14 0.66 0.14 1.345 0.08 1.345 0.08 0.73 0.06 0.73 0.06 0.6 0.08 0.6 0.08 0.54 0.14 0.54 0.14 0.6 0.49 0.6 0.49 0.54 0.55 0.54 0.55 0.6 0.9 0.6 0.9 0.54 0.96 0.54 0.96 0.6 1.31 0.6 1.31 0.54 1.37 0.54 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 0 1.77 0 1.65 0.285 1.65 0.285 0.9 0.345 0.9 0.345 1.65 0.695 1.65 0.695 0.9 0.755 0.9 0.755 1.65 1.105 1.65 1.105 0.9 1.165 0.9 1.165 1.65 1.515 1.65 1.515 1.225 1.575 1.225 1.575 1.65 2.045 1.65 2.045 0.975 2.105 0.975 2.105 1.65 2.455 1.65 2.455 1.245 2.515 1.245 2.515 1.65 2.835 1.65 2.835 1.275 2.955 1.275 2.955 1.335 2.895 1.335 2.895 1.65 4.365 1.65 4.365 1.54 4.485 1.54 4.485 1.65 4.69 1.65 4.69 1.37 4.63 1.37 4.63 1.31 4.75 1.31 4.75 1.65 5.53 1.65 5.53 1.24 5.59 1.24 5.59 1.65 6.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 5.59 0.06 5.59 0.44 5.53 0.44 5.53 0.06 4.725 0.06 4.725 0.29 4.785 0.29 4.785 0.35 4.665 0.35 4.665 0.06 4.085 0.06 4.085 0.17 3.965 0.17 3.965 0.06 2.515 0.06 2.515 0.45 2.455 0.45 2.455 0.06 2.105 0.06 2.105 0.52 2.045 0.52 2.045 0.06 1.605 0.06 1.605 0.2 1.545 0.2 1.545 0.06 1.165 0.06 1.165 0.485 1.105 0.485 1.105 0.06 0.755 0.06 0.755 0.485 0.695 0.485 0.695 0.06 0.345 0.06 0.345 0.485 0.285 0.485 0.285 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.795 0.465 5.75 0.465 5.75 0.6 5.37 0.6 5.37 1.08 5.795 1.08 5.795 1.265 5.735 1.265 5.735 1.14 5.37 1.14 5.37 1.33 5.03 1.33 5.03 1.37 4.91 1.37 4.91 1.21 4.265 1.21 4.265 1.37 3.9 1.37 3.9 1.31 4.205 1.31 4.205 1.15 4.97 1.15 4.97 1.27 5.31 1.27 5.31 0.685 5.25 0.685 5.25 0.54 5.69 0.54 5.69 0.405 5.735 0.405 5.735 0.345 5.795 0.345 ;
      POLYGON 5.15 1.17 5.09 1.17 5.09 0.83 4.535 0.83 4.535 0.77 5.09 0.77 5.09 0.345 5.15 0.345 ;
      POLYGON 4.99 0.635 4.93 0.635 4.93 0.51 4.505 0.51 4.505 0.35 4.245 0.35 4.245 0.89 3.885 0.89 3.885 0.99 3.945 0.99 3.945 1.05 3.825 1.05 3.825 0.515 3.57 0.515 3.57 0.395 3.63 0.395 3.63 0.455 3.885 0.455 3.885 0.83 4.185 0.83 4.185 0.29 4.565 0.29 4.565 0.45 4.99 0.45 ;
      POLYGON 4.83 0.67 4.405 0.67 4.405 0.93 4.485 0.93 4.485 1.05 4.105 1.05 4.105 1.21 3.7 1.21 3.7 1.235 3.64 1.235 3.64 0.955 3.665 0.955 3.665 0.675 3.41 0.675 3.41 0.505 3.35 0.505 3.35 0.445 3.47 0.445 3.47 0.615 3.725 0.615 3.725 1.15 4.045 1.15 4.045 0.99 4.345 0.99 4.345 0.45 4.405 0.45 4.405 0.61 4.83 0.61 ;
      POLYGON 3.565 0.855 3.2 0.855 3.2 0.64 3.28 0.64 3.28 0.775 3.565 0.775 ;
      POLYGON 3.495 1.235 3.435 1.235 3.435 1.015 2.425 1.015 2.425 0.88 2.365 0.88 2.365 0.82 2.485 0.82 2.485 0.955 3.04 0.955 3.04 0.445 3.25 0.445 3.25 0.505 3.1 0.505 3.1 0.955 3.495 0.955 ;
      POLYGON 3.29 1.235 3.23 1.235 3.23 1.175 2.72 1.175 2.72 1.235 2.66 1.235 2.66 1.115 3.29 1.115 ;
      POLYGON 2.76 0.695 2.265 0.695 2.265 0.975 2.31 0.975 2.31 1.365 2.25 1.365 2.25 1.035 2.205 1.035 2.205 0.695 1.9 0.695 1.9 1.095 1.84 1.095 1.84 0.76 1.53 0.76 1.53 0.82 1.47 0.82 1.47 0.7 1.84 0.7 1.84 0.54 1.9 0.54 1.9 0.635 2.25 0.635 2.25 0.47 2.31 0.47 2.31 0.635 2.7 0.635 2.7 0.575 2.76 0.575 ;
  END
END DFFSHQX8

MACRO DFFSRHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRHQX1 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6013 LAYER Metal1 ;
    ANTENNADIFFAREA 3.627875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2772 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.99170275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 102.24025975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.14 1.29 0.08 1.29 0.08 0.73 0.06 0.73 0.06 0.6 0.08 0.6 0.08 0.54 0.14 0.54 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.165 0.895 6.035 0.895 6.035 0.445 6.115 0.445 6.115 0.815 6.165 0.815 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.545 0.895 5.255 0.895 5.255 1.005 5.165 1.005 5.165 0.805 5.245 0.805 5.245 0.815 5.545 0.815 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 22.68608425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.99 1.44 3.68 1.44 3.68 1.28 3.36 1.28 3.36 1.345 2.295 1.345 2.295 1.2 1.9 1.2 1.9 1.26 1.46 1.26 1.46 0.835 1.42 0.835 1.42 0.775 1.54 0.775 1.54 0.92 1.52 0.92 1.52 1.2 1.84 1.2 1.84 1.14 2.355 1.14 2.355 1.285 3.3 1.285 3.3 1.22 3.74 1.22 3.74 1.38 3.99 1.38 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.32 0.895 1.035 0.895 1.035 0.79 0.925 0.79 0.925 0.71 1.115 0.71 1.115 0.815 1.32 0.815 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 1.77 0 1.77 0 1.65 0.285 1.65 0.285 1.08 0.345 1.08 0.345 1.65 1.14 1.65 1.14 1.215 1.08 1.215 1.08 1.155 1.2 1.155 1.2 1.65 2.075 1.65 2.075 1.3 2.195 1.3 2.195 1.36 2.135 1.36 2.135 1.65 3.52 1.65 3.52 1.44 3.46 1.44 3.46 1.38 3.58 1.38 3.58 1.65 4.44 1.65 4.44 1.31 4.38 1.31 4.38 1.25 4.5 1.25 4.5 1.65 5.27 1.65 5.27 1.265 5.33 1.265 5.33 1.65 6.11 1.65 6.11 0.995 6.17 0.995 6.17 1.65 6.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 0.06 6.275 0.06 6.275 0.635 6.215 0.635 6.215 0.06 5.33 0.06 5.33 0.48 5.27 0.48 5.27 0.06 4.295 0.06 4.295 0.48 4.235 0.48 4.235 0.06 1.285 0.06 1.285 0.45 1.225 0.45 1.225 0.06 0.345 0.06 0.345 0.575 0.285 0.575 0.285 0.06 0 0.06 0 -0.06 6.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.995 1.055 5.875 1.055 5.875 0.47 5.49 0.47 5.49 0.695 5.125 0.695 5.125 0.705 5.005 0.705 5.005 0.635 5.065 0.635 5.065 0.375 4.685 0.375 4.685 0.77 4.745 0.77 4.745 0.83 4.625 0.83 4.625 0.64 3.86 0.64 3.86 0.8 3.14 0.8 3.14 0.74 3.8 0.74 3.8 0.58 4.625 0.58 4.625 0.315 5.125 0.315 5.125 0.635 5.43 0.635 5.43 0.385 5.55 0.385 5.55 0.41 5.935 0.41 5.935 0.995 5.995 0.995 ;
      POLYGON 5.765 0.855 5.705 0.855 5.705 1.29 5.525 1.29 5.525 1.165 5.065 1.165 5.065 1.355 4.685 1.355 4.685 1.15 4.28 1.15 4.28 1.28 3.84 1.28 3.84 1.12 3.2 1.12 3.2 1.185 2.5 1.185 2.5 0.735 2.56 0.735 2.56 1.125 2.82 1.125 2.82 0.605 2.88 0.605 2.88 1.125 3.14 1.125 3.14 1.06 3.9 1.06 3.9 1.22 4.22 1.22 4.22 1.09 4.745 1.09 4.745 1.295 5.005 1.295 5.005 0.905 5.065 0.905 5.065 1.105 5.645 1.105 5.645 0.57 5.765 0.57 ;
      POLYGON 4.965 0.535 4.905 0.535 4.905 1.195 4.845 1.195 4.845 0.99 4.465 0.99 4.465 0.8 3.96 0.8 3.96 0.74 4.525 0.74 4.525 0.93 4.845 0.93 4.845 0.475 4.965 0.475 ;
      POLYGON 4.365 0.96 4.12 0.96 4.12 1.12 4 1.12 4 1.06 4.06 1.06 4.06 0.96 3.04 0.96 3.04 1.025 2.98 1.025 2.98 0.435 3.04 0.435 3.04 0.55 3.64 0.55 3.64 0.42 3.815 0.42 3.815 0.48 3.7 0.48 3.7 0.61 3.04 0.61 3.04 0.9 4.365 0.9 ;
      POLYGON 3.995 0.48 3.915 0.48 3.915 0.32 3.54 0.32 3.54 0.45 3.42 0.45 3.42 0.37 3.46 0.37 3.46 0.24 3.995 0.24 ;
      POLYGON 2.72 1.025 2.66 1.025 2.66 0.635 2.4 0.635 2.4 0.74 1.64 0.74 1.64 0.61 1.065 0.61 1.065 0.285 0.505 0.285 0.505 0.82 0.445 0.82 0.445 0.225 1.125 0.225 1.125 0.55 1.7 0.55 1.7 0.68 2.34 0.68 2.34 0.575 2.66 0.575 2.66 0.435 2.72 0.435 ;
      POLYGON 2.545 0.475 2.24 0.475 2.24 0.58 1.8 0.58 1.8 0.45 1.725 0.45 1.725 0.39 1.86 0.39 1.86 0.52 2.18 0.52 2.18 0.415 2.545 0.415 ;
      POLYGON 2.4 1.015 1.74 1.015 1.74 1.1 1.62 1.1 1.62 1.02 1.66 1.02 1.66 0.935 2.4 0.935 ;
      POLYGON 2.08 0.42 1.96 0.42 1.96 0.29 1.625 0.29 1.625 0.45 1.545 0.45 1.545 0.21 2.04 0.21 2.04 0.34 2.08 0.34 ;
      POLYGON 1.975 1.535 1.3 1.535 1.3 1.055 0.765 1.055 0.765 0.385 0.965 0.385 0.965 0.445 0.825 0.445 0.825 0.995 1.36 0.995 1.36 1.475 1.975 1.475 ;
      POLYGON 1.04 1.42 0.51 1.42 0.51 1.17 0.605 1.17 0.605 0.98 0.24 0.98 0.24 0.74 0.3 0.74 0.3 0.92 0.605 0.92 0.605 0.54 0.665 0.54 0.665 1.23 0.57 1.23 0.57 1.36 1.04 1.36 ;
  END
END DFFSRHQX1

MACRO DFFSRHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRHQX2 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6515 LAYER Metal1 ;
    ANTENNADIFFAREA 3.8552 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.30645 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.91548375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 93.92070475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.565 1.275 0.475 1.275 0.475 1.3 0.415 1.3 0.415 0.54 0.475 0.54 0.475 1.195 0.565 1.195 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.26 0.6 6.34 1.1 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.765 0.705 5.715 0.705 5.715 0.85 5.41 0.85 5.41 0.77 5.635 0.77 5.635 0.625 5.765 0.625 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 22.7184465 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.325 1.45 3.925 1.45 3.925 1.26 3.605 1.26 3.605 1.34 2.53 1.34 2.53 1.26 2.085 1.26 2.085 1.28 1.705 1.28 1.705 1.085 1.635 1.085 1.635 1.005 1.7 1.005 1.7 0.83 1.76 0.83 1.76 1.005 1.765 1.005 1.765 1.22 2.025 1.22 2.025 1.2 2.59 1.2 2.59 1.28 3.545 1.28 3.545 1.2 3.985 1.2 3.985 1.39 4.325 1.39 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.535 0.91 1.34 0.91 1.34 1.135 1.26 1.135 1.26 0.83 1.535 0.83 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 1.77 0 1.77 0 1.65 0.21 1.65 0.21 0.91 0.27 0.91 0.27 1.65 0.665 1.65 0.665 1.08 0.725 1.08 0.725 1.65 1.325 1.65 1.325 1.395 1.445 1.395 1.445 1.455 1.385 1.455 1.385 1.65 2.31 1.65 2.31 1.36 2.43 1.36 2.43 1.42 2.37 1.42 2.37 1.65 3.765 1.65 3.765 1.42 3.705 1.42 3.705 1.36 3.825 1.36 3.825 1.65 4.54 1.65 4.54 1.42 4.48 1.42 4.48 1.36 4.6 1.36 4.6 1.65 5.485 1.65 5.485 1.11 5.545 1.11 5.545 1.65 6.44 1.65 6.44 0.995 6.5 0.995 6.5 1.65 6.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 0.06 6.5 0.06 6.5 0.635 6.44 0.635 6.44 0.06 5.605 0.06 5.605 0.17 5.485 0.17 5.485 0.06 4.51 0.06 4.51 0.4 4.57 0.4 4.57 0.46 4.45 0.46 4.45 0.06 1.6 0.06 1.6 0.48 1.66 0.48 1.66 0.54 1.54 0.54 1.54 0.06 0.68 0.06 0.68 0.575 0.62 0.575 0.62 0.06 0.27 0.06 0.27 0.52 0.21 0.52 0.21 0.06 0 0.06 0 -0.06 6.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.16 1.02 6.1 1.02 6.1 0.435 5.385 0.435 5.385 0.67 5.31 0.67 5.31 0.745 5.25 0.745 5.25 0.61 5.325 0.61 5.325 0.35 4.93 0.35 4.93 0.855 4.99 0.855 4.99 0.915 4.87 0.915 4.87 0.62 4.105 0.62 4.105 0.78 3.385 0.78 3.385 0.72 4.045 0.72 4.045 0.56 4.87 0.56 4.87 0.29 5.385 0.29 5.385 0.375 6.16 0.375 ;
      POLYGON 5.985 0.63 5.925 0.63 5.925 1.01 5.75 1.01 5.75 1.135 5.69 1.135 5.69 1.01 5.31 1.01 5.31 1.295 4.93 1.295 4.93 1.26 4.085 1.26 4.085 1.1 3.445 1.1 3.445 1.18 2.745 1.18 2.745 0.83 2.685 0.83 2.685 0.77 2.805 0.77 2.805 1.12 3.065 1.12 3.065 0.61 3.125 0.61 3.125 1.12 3.385 1.12 3.385 1.04 4.145 1.04 4.145 1.2 4.99 1.2 4.99 1.235 5.25 1.235 5.25 0.845 5.31 0.845 5.31 0.95 5.865 0.95 5.865 0.57 5.985 0.57 ;
      POLYGON 5.225 0.51 5.15 0.51 5.15 1.135 5.09 1.135 5.09 1.075 4.71 1.075 4.71 0.78 4.205 0.78 4.205 0.72 4.77 0.72 4.77 1.015 5.09 1.015 5.09 0.45 5.225 0.45 ;
      POLYGON 4.61 0.94 4.365 0.94 4.365 1.1 4.245 1.1 4.245 1.04 4.305 1.04 4.305 0.94 3.285 0.94 3.285 1.02 3.225 1.02 3.225 0.51 3.11 0.51 3.11 0.39 3.17 0.39 3.17 0.45 3.285 0.45 3.285 0.56 3.825 0.56 3.825 0.485 3.945 0.485 3.945 0.545 3.885 0.545 3.885 0.62 3.285 0.62 3.285 0.88 4.61 0.88 ;
      POLYGON 4.285 0.46 4.045 0.46 4.045 0.385 3.725 0.385 3.725 0.46 3.605 0.46 3.605 0.38 3.645 0.38 3.645 0.305 4.125 0.305 4.125 0.38 4.285 0.38 ;
      POLYGON 2.965 1.02 2.905 1.02 2.905 0.67 2.585 0.67 2.585 0.89 1.865 0.89 1.865 0.73 1.31 0.73 1.31 0.435 0.84 0.435 0.84 0.82 0.78 0.82 0.78 0.375 1.37 0.375 1.37 0.67 1.925 0.67 1.925 0.83 2.525 0.83 2.525 0.61 2.905 0.61 2.905 0.45 2.965 0.45 ;
      POLYGON 2.79 0.51 2.425 0.51 2.425 0.73 2.025 0.73 2.025 0.57 1.95 0.57 1.95 0.51 2.085 0.51 2.085 0.67 2.365 0.67 2.365 0.45 2.79 0.45 ;
      POLYGON 2.645 1.05 1.925 1.05 1.925 1.12 1.865 1.12 1.865 0.99 2.645 0.99 ;
      POLYGON 2.265 0.57 2.185 0.57 2.185 0.41 1.85 0.41 1.85 0.57 1.77 0.57 1.77 0.33 2.265 0.33 ;
      POLYGON 2.21 1.525 1.545 1.525 1.545 1.295 1.1 1.295 1.1 0.595 1.15 0.595 1.15 0.535 1.21 0.535 1.21 0.655 1.16 0.655 1.16 1.235 1.605 1.235 1.605 1.465 2.21 1.465 ;
      POLYGON 1.225 1.55 0.87 1.55 0.87 1.18 0.94 1.18 0.94 0.98 0.575 0.98 0.575 0.74 0.635 0.74 0.635 0.92 0.94 0.92 0.94 0.54 1 0.54 1 1.24 0.93 1.24 0.93 1.49 1.225 1.49 ;
  END
END DFFSRHQX2

MACRO DFFSRHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRHQX4 0 0 ;
  SIZE 7.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 18.28478975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.205 1.34 4.545 1.34 4.545 1.285 4.225 1.285 4.225 1.405 3.365 1.405 3.365 1.065 3.165 1.065 3.165 1.085 3.035 1.085 3.035 1.065 2.975 1.065 2.975 1.005 3.425 1.005 3.425 1.345 4.165 1.345 4.165 1.225 4.605 1.225 4.605 1.28 5.205 1.28 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.37 0.745 7.085 0.745 7.085 0.84 7.005 0.84 7.005 0.625 7.37 0.625 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.695793 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.275 0.815 6.585 0.945 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.605 0.625 1.775 0.865 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.06285 LAYER Metal1 ;
    ANTENNADIFFAREA 4.4279 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.388125 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.4678905 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 82.00966175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.905 1.34 0.845 1.34 0.845 0.73 0.495 0.73 0.495 1.34 0.435 1.34 0.435 0.415 0.495 0.415 0.495 0.6 0.54 0.6 0.54 0.67 0.845 0.67 0.845 0.415 0.905 0.415 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.4 1.77 0 1.77 0 1.65 0.23 1.65 0.23 0.95 0.29 0.95 0.29 1.65 0.64 1.65 0.64 0.95 0.7 0.95 0.7 1.65 1.075 1.65 1.075 1.03 1.135 1.03 1.135 1.65 1.485 1.65 1.485 1.125 1.545 1.125 1.545 1.65 2.245 1.65 2.245 1.47 2.185 1.47 2.185 1.41 2.305 1.41 2.305 1.65 2.89 1.65 2.89 1.54 3.01 1.54 3.01 1.65 4.385 1.65 4.385 1.445 4.325 1.445 4.325 1.385 4.445 1.385 4.445 1.65 5.33 1.65 5.33 1.25 5.45 1.25 5.45 1.31 5.39 1.31 5.39 1.65 6.35 1.65 6.35 1.25 6.41 1.25 6.41 1.65 7.17 1.65 7.17 0.995 7.23 0.995 7.23 1.65 7.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.4 0.06 7.175 0.06 7.175 0.525 7.115 0.525 7.115 0.06 6.335 0.06 6.335 0.55 6.275 0.55 6.275 0.06 5.52 0.06 5.52 0.455 5.46 0.455 5.46 0.06 3.155 0.06 3.155 0.17 3.035 0.17 3.035 0.06 1.575 0.06 1.575 0.365 1.455 0.365 1.455 0.305 1.515 0.305 1.515 0.06 1.11 0.06 1.11 0.395 1.05 0.395 1.05 0.06 0.7 0.06 0.7 0.395 0.64 0.395 0.64 0.06 0.29 0.06 0.29 0.395 0.23 0.395 0.23 0.06 0 0.06 0 -0.06 7.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.965 1 6.845 1 6.845 0.385 6.495 0.385 6.495 0.655 6.555 0.655 6.555 0.715 6.015 0.715 6.015 1.34 5.575 1.34 5.575 1.15 4.705 1.15 4.705 1.125 4.065 1.125 4.065 1.245 3.685 1.245 3.685 0.745 3.745 0.745 3.745 0.415 3.425 0.415 3.425 0.745 3.305 0.745 3.305 0.685 3.365 0.685 3.365 0.355 3.805 0.355 3.805 0.805 3.745 0.805 3.745 1.185 4.005 1.185 4.005 1.065 4.765 1.065 4.765 1.09 5.575 1.09 5.575 0.93 5.695 0.93 5.695 0.99 5.635 0.99 5.635 1.28 5.955 1.28 5.955 0.655 6.435 0.655 6.435 0.325 6.905 0.325 6.905 0.94 6.965 0.94 ;
      POLYGON 6.745 1.105 6.615 1.105 6.615 1.275 6.555 1.275 6.555 1.105 6.115 1.105 6.115 0.89 6.175 0.89 6.175 1.045 6.685 1.045 6.685 0.545 6.595 0.545 6.595 0.485 6.745 0.485 ;
      POLYGON 5.855 1.18 5.795 1.18 5.795 0.555 5.68 0.555 5.68 0.67 5.185 0.67 5.185 0.61 5.62 0.61 5.62 0.495 5.795 0.495 5.795 0.42 5.855 0.42 ;
      POLYGON 5.695 0.83 5.025 0.83 5.025 0.795 4.065 0.795 4.065 0.735 5.085 0.735 5.085 0.77 5.695 0.77 ;
      POLYGON 5.475 0.99 4.865 0.99 4.865 0.965 3.905 0.965 3.905 1.085 3.845 1.085 3.845 0.905 3.905 0.905 3.905 0.485 3.965 0.485 3.965 0.575 4.85 0.575 4.85 0.5 4.97 0.5 4.97 0.56 4.91 0.56 4.91 0.635 3.965 0.635 3.965 0.905 4.925 0.905 4.925 0.93 5.475 0.93 ;
      POLYGON 5.15 0.505 5.07 0.505 5.07 0.4 4.75 0.4 4.75 0.475 4.63 0.475 4.63 0.395 4.67 0.395 4.67 0.32 5.15 0.32 ;
      POLYGON 3.645 0.575 3.585 0.575 3.585 1.245 3.525 1.245 3.525 0.905 2.875 0.905 2.875 1.045 2.365 1.045 2.365 1.31 1.645 1.31 1.645 1.025 1.44 1.025 1.44 0.87 1.5 0.87 1.5 0.965 1.705 0.965 1.705 1.25 2.305 1.25 2.305 0.985 2.815 0.985 2.815 0.845 3.525 0.845 3.525 0.515 3.645 0.515 ;
      POLYGON 3.265 0.575 2.875 0.575 2.875 0.405 2.555 0.405 2.555 0.48 2.435 0.48 2.435 0.42 2.495 0.42 2.495 0.345 2.935 0.345 2.935 0.515 3.265 0.515 ;
      POLYGON 3.265 1.265 2.685 1.265 2.685 1.145 2.765 1.145 2.765 1.185 3.265 1.185 ;
      POLYGON 3.265 1.55 3.145 1.55 3.145 1.44 2.525 1.44 2.525 1.47 2.405 1.47 2.405 1.41 2.465 1.41 2.465 1.38 3.205 1.38 3.205 1.49 3.265 1.49 ;
      POLYGON 2.775 0.565 2.715 0.565 2.715 0.885 2.115 0.885 2.115 0.565 2.055 0.565 2.055 0.505 2.175 0.505 2.175 0.825 2.655 0.825 2.655 0.505 2.775 0.505 ;
      POLYGON 2.555 0.725 2.275 0.725 2.275 0.345 1.735 0.345 1.735 0.525 1.34 0.525 1.34 1.15 1.28 1.15 1.28 0.665 1.005 0.665 1.005 0.605 1.28 0.605 1.28 0.36 1.34 0.36 1.34 0.465 1.675 0.465 1.675 0.285 2.335 0.285 2.335 0.665 2.555 0.665 ;
      POLYGON 2.015 0.83 1.955 0.83 1.955 1.11 1.885 1.11 1.885 1.15 1.805 1.15 1.805 1.03 1.875 1.03 1.875 0.525 1.835 0.525 1.835 0.445 1.955 0.445 1.955 0.75 2.015 0.75 ;
  END
END DFFSRHQX4

MACRO DFFSRHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRHQX8 0 0 ;
  SIZE 7.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.46 0.655 7.54 1.155 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.975 0.705 6.885 0.705 6.885 0.865 6.765 0.865 6.765 0.625 6.835 0.625 6.835 0.495 6.975 0.495 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 22.459547 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.59 1.44 5.28 1.44 5.28 1.28 4.96 1.28 4.96 1.345 3.9 1.345 3.9 1.185 3.48 1.185 3.48 1.265 3.08 1.265 3.08 0.92 3.06 0.92 3.06 0.79 3.14 0.79 3.14 1.205 3.42 1.205 3.42 1.125 3.96 1.125 3.96 1.285 4.9 1.285 4.9 1.22 5.34 1.22 5.34 1.38 5.59 1.38 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.66 0.6 2.74 1.1 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4053 LAYER Metal1 ;
    ANTENNADIFFAREA 4.94025 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.545625 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.07386025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 63.53814425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.37 0.65 1.325 0.65 1.325 0.9 1.37 0.9 1.37 1.345 1.31 1.345 1.31 0.96 1.265 0.96 1.265 0.8 0.96 0.8 0.96 1.345 0.9 1.345 0.9 0.705 0.55 0.705 0.55 1.345 0.49 1.345 0.49 0.705 0.14 0.705 0.14 1.345 0.08 1.345 0.08 0.73 0.06 0.73 0.06 0.6 0.08 0.6 0.08 0.54 0.14 0.54 0.14 0.645 0.49 0.645 0.49 0.54 0.55 0.54 0.55 0.645 0.9 0.645 0.9 0.54 0.96 0.54 0.96 0.74 1.265 0.74 1.265 0.59 1.31 0.59 1.31 0.53 1.37 0.53 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.8 1.77 0 1.77 0 1.65 0.285 1.65 0.285 0.9 0.345 0.9 0.345 1.65 0.695 1.65 0.695 0.9 0.755 0.9 0.755 1.65 1.105 1.65 1.105 0.9 1.165 0.9 1.165 1.65 1.515 1.65 1.515 0.955 1.575 0.955 1.575 1.65 1.925 1.65 1.925 1.08 1.985 1.08 1.985 1.65 2.76 1.65 2.76 1.42 2.7 1.42 2.7 1.36 2.82 1.36 2.82 1.65 3.68 1.65 3.68 1.285 3.8 1.285 3.8 1.345 3.74 1.345 3.74 1.65 5.12 1.65 5.12 1.44 5.06 1.44 5.06 1.38 5.18 1.38 5.18 1.65 6.04 1.65 6.04 1.31 5.98 1.31 5.98 1.25 6.1 1.25 6.1 1.65 6.84 1.65 6.84 1.125 6.9 1.125 6.9 1.65 7.525 1.65 7.525 1.255 7.585 1.255 7.585 1.65 7.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.8 0.06 7.62 0.06 7.62 0.2 7.56 0.2 7.56 0.06 6.96 0.06 6.96 0.17 6.84 0.17 6.84 0.06 5.895 0.06 5.895 0.48 5.835 0.48 5.835 0.06 3.01 0.06 3.01 0.17 2.89 0.17 2.89 0.06 1.985 0.06 1.985 0.52 1.925 0.52 1.925 0.06 1.575 0.06 1.575 0.52 1.515 0.52 1.515 0.06 1.165 0.06 1.165 0.485 1.105 0.485 1.105 0.06 0.755 0.06 0.755 0.485 0.695 0.485 0.695 0.06 0.345 0.06 0.345 0.485 0.285 0.485 0.285 0.06 0 0.06 0 -0.06 7.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.455 0.555 7.36 0.555 7.36 1.28 7.3 1.28 7.3 0.495 7.395 0.495 7.395 0.395 6.665 0.395 6.665 0.735 6.605 0.735 6.605 0.375 6.285 0.375 6.285 0.77 6.345 0.77 6.345 0.83 6.225 0.83 6.225 0.64 5.46 0.64 5.46 0.8 4.74 0.8 4.74 0.74 5.4 0.74 5.4 0.58 6.225 0.58 6.225 0.315 6.665 0.315 6.665 0.335 7.455 0.335 ;
      POLYGON 7.195 0.58 7.135 0.58 7.135 1.025 7.105 1.025 7.105 1.15 7.045 1.15 7.045 1.025 6.665 1.025 6.665 1.31 6.285 1.31 6.285 1.15 5.88 1.15 5.88 1.28 5.44 1.28 5.44 1.12 4.8 1.12 4.8 1.185 4.1 1.185 4.1 0.745 4.16 0.745 4.16 1.125 4.42 1.125 4.42 0.605 4.48 0.605 4.48 1.125 4.74 1.125 4.74 1.06 5.5 1.06 5.5 1.22 5.82 1.22 5.82 1.09 6.345 1.09 6.345 1.25 6.605 1.25 6.605 0.86 6.665 0.86 6.665 0.965 7.075 0.965 7.075 0.52 7.195 0.52 ;
      POLYGON 6.505 1.15 6.445 1.15 6.445 0.99 6.065 0.99 6.065 0.8 5.56 0.8 5.56 0.74 6.125 0.74 6.125 0.93 6.445 0.93 6.445 0.535 6.385 0.535 6.385 0.475 6.505 0.475 ;
      POLYGON 5.965 0.96 5.72 0.96 5.72 1.12 5.6 1.12 5.6 1.06 5.66 1.06 5.66 0.96 4.64 0.96 4.64 1.025 4.58 1.025 4.58 0.435 4.64 0.435 4.64 0.55 5.24 0.55 5.24 0.42 5.415 0.42 5.415 0.48 5.3 0.48 5.3 0.61 4.64 0.61 4.64 0.9 5.965 0.9 ;
      POLYGON 5.595 0.48 5.515 0.48 5.515 0.32 5.14 0.32 5.14 0.45 5.02 0.45 5.02 0.37 5.06 0.37 5.06 0.24 5.595 0.24 ;
      POLYGON 4.405 0.505 4.32 0.505 4.32 1.025 4.26 1.025 4.26 0.645 4 0.645 4 0.76 3.24 0.76 3.24 0.685 2.99 0.685 2.99 0.34 2.145 0.34 2.145 0.82 2.085 0.82 2.085 0.28 3.05 0.28 3.05 0.625 3.3 0.625 3.3 0.7 3.94 0.7 3.94 0.585 4.26 0.585 4.26 0.445 4.345 0.445 4.345 0.385 4.405 0.385 ;
      POLYGON 4.16 0.485 3.84 0.485 3.84 0.6 3.4 0.6 3.4 0.525 3.33 0.525 3.33 0.465 3.46 0.465 3.46 0.54 3.78 0.54 3.78 0.425 4.16 0.425 ;
      POLYGON 4 1.025 3.32 1.025 3.32 1.105 3.24 1.105 3.24 0.945 3.92 0.945 3.92 0.905 4 0.905 ;
      POLYGON 3.68 0.44 3.56 0.44 3.56 0.365 3.23 0.365 3.23 0.47 3.15 0.47 3.15 0.285 3.64 0.285 3.64 0.36 3.68 0.36 ;
      POLYGON 3.58 1.535 2.92 1.535 2.92 1.26 2.495 1.26 2.495 0.44 2.685 0.44 2.685 0.5 2.555 0.5 2.555 1.2 2.98 1.2 2.98 1.475 3.58 1.475 ;
      POLYGON 2.65 1.55 2.13 1.55 2.13 1.225 2.245 1.225 2.245 0.98 1.78 0.98 1.78 1.345 1.72 1.345 1.72 0.805 1.425 0.805 1.425 0.745 1.72 0.745 1.72 0.54 1.78 0.54 1.78 0.92 2.245 0.92 2.245 0.54 2.305 0.54 2.305 1.285 2.19 1.285 2.19 1.49 2.65 1.49 ;
  END
END DFFSRHQX8

MACRO DFFSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRX1 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.50855 LAYER Metal1 ;
    ANTENNADIFFAREA 3.64745 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2529 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.87327 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 106.049822 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.09 1.17 1.03 1.17 1.03 1.11 0.86 1.11 0.86 0.98 0.88 0.98 0.88 0.4 1.02 0.4 1.02 0.34 1.08 0.34 1.08 0.46 0.94 0.46 0.94 1.05 1.09 1.05 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.50855 LAYER Metal1 ;
    ANTENNADIFFAREA 3.64745 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2529 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.87327 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 106.049822 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.325 1.29 0.245 1.29 0.245 0.73 0.06 0.73 0.06 0.6 0.245 0.6 0.245 0.54 0.325 0.54 ;
    END
  END QN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.54 0.54 6.48 0.54 6.48 0.85 6.4 0.85 6.4 0.46 6.46 0.46 6.46 0.41 6.54 0.41 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.94 0.925 5.86 0.925 5.86 0.87 5.68 0.87 5.68 0.605 5.76 0.605 5.76 0.79 5.94 0.79 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 35.04629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.855 0.92 3.945 0.92 3.945 0.36 3.365 0.36 3.365 0.865 2.265 0.865 2.265 0.805 3.305 0.805 3.305 0.705 3.235 0.705 3.235 0.625 3.305 0.625 3.305 0.3 4.005 0.3 4.005 0.86 4.855 0.86 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.445 0.8 1.365 0.8 1.365 0.895 1.04 0.895 1.04 0.815 1.285 0.815 1.285 0.72 1.445 0.72 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 1.77 0 1.77 0 1.65 0.5 1.65 0.5 1.285 0.56 1.285 0.56 1.65 1.235 1.65 1.235 0.995 1.295 0.995 1.295 1.65 2.135 1.65 2.135 1.38 2.195 1.38 2.195 1.65 2.92 1.65 2.92 1.305 2.98 1.305 2.98 1.65 4.13 1.65 4.13 1.54 4.25 1.54 4.25 1.65 4.905 1.65 4.905 1.54 5.025 1.54 5.025 1.65 5.84 1.65 5.84 1.51 5.9 1.51 5.9 1.65 6.445 1.65 6.445 1.29 6.505 1.29 6.505 1.65 6.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 0.06 6.465 0.06 6.465 0.2 6.405 0.2 6.405 0.06 5.77 0.06 5.77 0.505 5.71 0.505 5.71 0.06 5.025 0.06 5.025 0.17 4.905 0.17 4.905 0.06 2.255 0.06 2.255 0.495 2.135 0.495 2.135 0.435 2.195 0.435 2.195 0.06 1.285 0.06 1.285 0.445 1.225 0.445 1.225 0.06 0.56 0.06 0.56 0.2 0.5 0.2 0.5 0.06 0 0.06 0 -0.06 6.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.3 1.315 6.24 1.315 6.24 1.245 5.74 1.245 5.74 1.43 4.35 1.43 4.35 1.4 3.7 1.4 3.7 1.34 4.41 1.34 4.41 1.37 5.68 1.37 5.68 1.185 6.24 1.185 6.24 0.54 6.3 0.54 ;
      POLYGON 6.1 1.085 5.58 1.085 5.58 1.27 4.51 1.27 4.51 1.24 3.6 1.24 3.6 1.365 3.285 1.365 3.285 1.305 3.54 1.305 3.54 1.18 3.625 1.18 3.625 0.8 3.685 0.8 3.685 1.18 4.57 1.18 4.57 1.21 5.14 1.21 5.14 0.73 5.2 0.73 5.2 1.21 5.52 1.21 5.52 0.83 5.58 0.83 5.58 1.025 6.04 1.025 6.04 0.535 6.1 0.535 ;
      POLYGON 5.42 1.11 5.3 1.11 5.3 0.63 5.205 0.63 5.205 0.44 4.63 0.44 4.63 0.38 5.265 0.38 5.265 0.57 5.36 0.57 5.36 1.05 5.42 1.05 ;
      POLYGON 5.03 0.825 5.015 0.825 5.015 1.08 3.785 1.08 3.785 0.46 3.845 0.46 3.845 1.02 4.955 1.02 4.955 0.76 4.31 0.76 4.31 0.535 4.37 0.535 4.37 0.7 5.03 0.7 ;
      POLYGON 4.79 0.6 4.47 0.6 4.47 0.435 4.165 0.435 4.165 0.63 4.105 0.63 4.105 0.375 4.53 0.375 4.53 0.54 4.79 0.54 ;
      POLYGON 3.525 1.025 3.44 1.025 3.44 1.12 3.38 1.12 3.38 1.025 2.1 1.025 2.1 0.815 2.16 0.815 2.16 0.965 3.465 0.965 3.465 0.46 3.525 0.46 ;
      RECT 2.455 1.125 3.265 1.205 ;
      POLYGON 3.205 0.525 3.135 0.525 3.135 0.705 2.715 0.705 2.715 0.55 2.69 0.55 2.69 0.43 2.77 0.43 2.77 0.485 2.795 0.485 2.795 0.625 3.055 0.625 3.055 0.445 3.205 0.445 ;
      POLYGON 2.955 0.525 2.895 0.525 2.895 0.33 2.545 0.33 2.545 0.525 2.485 0.525 2.485 0.27 2.955 0.27 ;
      POLYGON 2.82 1.365 2.295 1.365 2.295 1.28 1.465 1.28 1.465 0.9 1.545 0.9 1.545 0.465 1.605 0.465 1.605 0.96 1.525 0.96 1.525 1.22 2.355 1.22 2.355 1.305 2.82 1.305 ;
      POLYGON 2.615 0.69 1.875 0.69 1.875 1.12 1.815 1.12 1.815 0.63 1.94 0.63 1.94 0.365 1.445 0.365 1.445 0.62 1.185 0.62 1.185 0.715 1.065 0.715 1.065 0.56 1.385 0.56 1.385 0.305 2 0.305 2 0.63 2.615 0.63 ;
      POLYGON 0.76 1.02 0.68 1.02 0.68 0.79 0.425 0.79 0.425 0.71 0.68 0.71 0.68 0.54 0.76 0.54 ;
  END
END DFFSRX1

MACRO DFFSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRX2 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.237025 LAYER Metal1 ;
    ANTENNADIFFAREA 4.336925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318375 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.30828425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 102.492344 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.455 0.65 7.34 0.65 7.34 0.915 7.365 0.915 7.365 1.305 7.285 1.305 7.285 1.11 7.26 1.11 7.26 0.57 7.455 0.57 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.237025 LAYER Metal1 ;
    ANTENNADIFFAREA 4.336925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.318375 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.30828425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 102.492344 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.96 1.305 6.88 1.305 6.88 1.11 6.86 1.11 6.86 0.98 6.88 0.98 6.88 0.54 6.96 0.54 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.62 1.085 6.42 1.085 6.42 1.005 6.54 1.005 6.54 0.705 6.62 0.705 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2322 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.16666675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 76.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.835 0.815 1.995 1.065 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.02 1.03 0.655 1.03 0.655 0.815 0.965 0.815 0.965 0.95 1.02 0.95 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.235 0.815 0.155 0.815 0.155 0.54 0.06 0.54 0.06 0.41 0.14 0.41 0.14 0.46 0.235 0.46 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 1.77 0 1.77 0 1.65 0.17 1.65 0.17 1.285 0.23 1.285 0.23 1.65 0.77 1.65 0.77 1.29 0.83 1.29 0.83 1.65 1.78 1.65 1.78 1.51 1.84 1.51 1.84 1.65 2.635 1.65 2.635 1.415 2.755 1.415 2.755 1.475 2.695 1.475 2.695 1.65 4.02 1.65 4.02 1.415 4.14 1.415 4.14 1.475 4.08 1.475 4.08 1.65 5.66 1.65 5.66 1.55 5.6 1.55 5.6 1.49 5.72 1.49 5.72 1.65 6.69 1.65 6.69 1.185 6.75 1.185 6.75 1.65 7.1 1.65 7.1 0.93 7.16 0.93 7.16 1.65 7.51 1.65 7.51 1.01 7.57 1.01 7.57 1.65 8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 0.06 7.72 0.06 7.72 0.17 7.6 0.17 7.6 0.06 7.22 0.06 7.22 0.17 7.1 0.17 7.1 0.06 6.75 0.06 6.75 0.17 6.63 0.17 6.63 0.06 5.775 0.06 5.775 0.54 5.715 0.54 5.715 0.06 1.78 0.06 1.78 0.495 1.84 0.495 1.84 0.555 1.72 0.555 1.72 0.06 0.955 0.06 0.955 0.2 0.895 0.2 0.895 0.06 0.23 0.06 0.23 0.2 0.17 0.2 0.17 0.06 0 0.06 0 -0.06 8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.885 0.63 7.775 0.63 7.775 1.035 7.715 1.035 7.715 0.815 7.44 0.815 7.44 0.755 7.715 0.755 7.715 0.57 7.885 0.57 ;
      POLYGON 7.88 0.44 7.12 0.44 7.12 0.83 7.06 0.83 7.06 0.44 6.78 0.44 6.78 0.83 6.72 0.83 6.72 0.44 6.04 0.44 6.04 1.245 5.98 1.245 5.98 0.705 5.42 0.705 5.42 0.645 5.98 0.645 5.98 0.38 7.76 0.38 7.76 0.375 7.88 0.375 ;
      POLYGON 6.575 0.605 6.32 0.605 6.32 1.185 6.545 1.185 6.545 1.405 5.82 1.405 5.82 1.185 4.4 1.185 4.4 1.155 3.915 1.155 3.915 1.095 4.46 1.095 4.46 1.125 5.88 1.125 5.88 1.345 6.485 1.345 6.485 1.245 6.26 1.245 6.26 0.545 6.575 0.545 ;
      POLYGON 5.88 0.865 4.72 0.865 4.72 0.835 3.555 0.835 3.555 1.02 3.495 1.02 3.495 0.43 3.555 0.43 3.555 0.775 4.78 0.775 4.78 0.805 5.88 0.805 ;
      POLYGON 5.6 0.51 5.48 0.51 5.48 0.375 5.16 0.375 5.16 0.51 5.04 0.51 5.04 0.43 5.08 0.43 5.08 0.295 5.56 0.295 5.56 0.43 5.6 0.43 ;
      POLYGON 5.5 1.345 4.24 1.345 4.24 1.315 3.555 1.315 3.555 1.34 2.855 1.34 2.855 1.315 2.535 1.315 2.535 1.545 1.94 1.545 1.94 1.485 2.475 1.485 2.475 1.255 2.915 1.255 2.915 1.28 3.495 1.28 3.495 1.255 4.3 1.255 4.3 1.285 5.5 1.285 ;
      POLYGON 5.47 1.025 4.56 1.025 4.56 0.995 3.76 0.995 3.76 1.055 3.7 1.055 3.7 0.935 4.62 0.935 4.62 0.965 5.47 0.965 ;
      POLYGON 5.38 0.535 5.32 0.535 5.32 0.67 4.88 0.67 4.88 0.52 3.67 0.52 3.67 0.46 4.94 0.46 4.94 0.61 5.26 0.61 5.26 0.475 5.38 0.475 ;
      POLYGON 3.635 0.22 3.395 0.22 3.395 1.18 3.015 1.18 3.015 1.155 2.375 1.155 2.375 1.385 1.68 1.385 1.68 1.475 1.28 1.475 1.28 0.77 1.22 0.77 1.22 0.715 0.675 0.715 0.675 0.655 0.735 0.655 0.735 0.335 0.395 0.335 0.395 1.02 0.335 1.02 0.335 0.275 0.795 0.275 0.795 0.655 1.28 0.655 1.28 0.71 1.34 0.71 1.34 1.415 1.62 1.415 1.62 1.325 2.315 1.325 2.315 1.095 3.075 1.095 3.075 1.12 3.335 1.12 3.335 0.16 3.635 0.16 ;
      POLYGON 3.235 1.02 3.175 1.02 3.175 0.96 2.155 0.96 2.155 1.165 2.215 1.165 2.215 1.225 1.675 1.225 1.675 0.96 1.735 0.96 1.735 1.165 2.095 1.165 2.095 0.9 2.38 0.9 2.38 0.61 2.36 0.61 2.36 0.49 2.42 0.49 2.42 0.56 2.44 0.56 2.44 0.9 3.175 0.9 3.175 0.43 3.235 0.43 ;
      POLYGON 2.625 0.585 2.565 0.585 2.565 0.39 2.215 0.39 2.215 0.555 2.095 0.555 2.095 0.495 2.155 0.495 2.155 0.33 2.625 0.33 ;
      POLYGON 2.28 0.74 2.16 0.74 2.16 0.715 1.5 0.715 1.5 1.315 1.44 1.315 1.44 0.49 1.5 0.49 1.5 0.655 2.22 0.655 2.22 0.68 2.28 0.68 ;
      POLYGON 1.18 1.19 0.625 1.19 0.625 1.315 0.495 1.315 0.495 0.495 0.575 0.495 0.575 0.435 0.635 0.435 0.635 0.555 0.555 0.555 0.555 1.13 1.12 1.13 1.12 1.025 1.18 1.025 ;
  END
END DFFSRX2

MACRO DFFSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRX4 0 0 ;
  SIZE 8.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7 LAYER Metal1 ;
    ANTENNADIFFAREA 4.921675 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4716 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.966073 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 78.816794 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.545 0.51 7.14 0.51 7.14 0.915 7.485 0.915 7.485 1.305 7.425 1.305 7.425 0.975 7.045 0.975 7.045 1.305 6.985 1.305 6.985 0.915 7.06 0.915 7.06 0.51 6.955 0.51 6.955 0.45 7.545 0.45 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.7 LAYER Metal1 ;
    ANTENNADIFFAREA 4.921675 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4716 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.966073 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 78.816794 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.605 0.5 6.14 0.5 6.14 0.915 6.555 0.915 6.555 1.305 6.495 1.305 6.495 0.975 6.12 0.975 6.12 1.305 6.06 1.305 6.06 0.6 6.08 0.6 6.08 0.5 6.015 0.5 6.015 0.44 6.605 0.44 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.51 0.895 3.195 0.895 3.195 0.815 3.235 0.815 3.235 0.63 3.51 0.63 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.095 0.895 2.78 0.895 2.78 0.815 2.835 0.815 2.835 0.63 3.095 0.63 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.765 1.085 0.445 1.085 0.445 1.005 0.58 1.005 0.58 0.825 0.765 0.825 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.63 0.34 1.13 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.2 1.77 0 1.77 0 1.65 0.42 1.65 0.42 1.23 0.48 1.23 0.48 1.65 1.43 1.65 1.43 1.49 1.55 1.49 1.55 1.55 1.49 1.55 1.49 1.65 1.86 1.65 1.86 1.55 1.8 1.55 1.8 1.49 1.92 1.49 1.92 1.65 3.13 1.65 3.13 1.375 3.07 1.375 3.07 1.315 3.19 1.315 3.19 1.65 4.785 1.65 4.785 1.185 4.845 1.185 4.845 1.65 5.3 1.65 5.3 1.185 5.36 1.185 5.36 1.65 5.75 1.65 5.75 0.995 5.81 0.995 5.81 1.65 6.265 1.65 6.265 1.075 6.325 1.075 6.325 1.65 6.72 1.65 6.72 0.915 6.78 0.915 6.78 1.65 7.22 1.65 7.22 1.075 7.28 1.075 7.28 1.65 7.655 1.65 7.655 0.955 7.715 0.955 7.715 1.65 8.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.2 0.06 7.865 0.06 7.865 0.4 7.805 0.4 7.805 0.06 7.31 0.06 7.31 0.17 7.19 0.17 7.19 0.06 6.84 0.06 6.84 0.17 6.72 0.17 6.72 0.06 6.37 0.06 6.37 0.17 6.25 0.17 6.25 0.06 5.695 0.06 5.695 0.365 5.755 0.365 5.755 0.425 5.635 0.425 5.635 0.06 5.315 0.06 5.315 0.455 5.255 0.455 5.255 0.06 3.265 0.06 3.265 0.37 3.145 0.37 3.145 0.31 3.205 0.31 3.205 0.06 1.555 0.06 1.555 0.17 1.435 0.17 1.435 0.06 0.5 0.06 0.5 0.2 0.44 0.2 0.44 0.06 0 0.06 0 -0.06 8.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 8.07 0.54 8.045 0.54 8.045 0.855 7.92 0.855 7.92 1.305 7.86 1.305 7.86 0.855 7.585 0.855 7.585 0.785 7.705 0.785 7.705 0.795 7.985 0.795 7.985 0.48 8.01 0.48 8.01 0.42 8.07 0.42 ;
      POLYGON 7.885 0.695 7.765 0.695 7.765 0.685 7.645 0.685 7.645 0.34 5.915 0.34 5.915 0.645 5.605 0.645 5.605 0.785 5.96 0.785 5.96 0.845 5.605 0.845 5.605 1.305 5.545 1.305 5.545 0.645 4.99 0.645 4.99 0.585 5.46 0.585 5.46 0.42 5.52 0.42 5.52 0.585 5.855 0.585 5.855 0.28 7.705 0.28 7.705 0.625 7.825 0.625 7.825 0.635 7.885 0.635 ;
      POLYGON 5.445 0.925 4.15 0.925 4.15 1.145 4.09 1.145 4.09 0.63 4.06 0.63 4.06 0.51 4.12 0.51 4.12 0.57 4.15 0.57 4.15 0.865 5.385 0.865 5.385 0.805 5.445 0.805 ;
      POLYGON 5.185 1.18 5.065 1.18 5.065 1.085 4.265 1.085 4.265 1.025 5.125 1.025 5.125 1.12 5.185 1.12 ;
      POLYGON 5.11 0.455 5.05 0.455 5.05 0.26 4.71 0.26 4.71 0.425 4.59 0.425 4.59 0.365 4.65 0.365 4.65 0.2 5.11 0.2 ;
      POLYGON 4.89 0.605 4.41 0.605 4.41 0.485 4.49 0.485 4.49 0.525 4.81 0.525 4.81 0.36 4.89 0.36 ;
      POLYGON 4.79 0.765 4.25 0.765 4.25 0.37 3.47 0.37 3.47 0.47 3.67 0.47 3.67 1.02 3.61 1.02 3.61 0.53 2.985 0.53 2.985 0.31 2.55 0.31 2.55 0.25 3.045 0.25 3.045 0.47 3.41 0.47 3.41 0.31 4.31 0.31 4.31 0.705 4.79 0.705 ;
      POLYGON 4.245 1.4 3.29 1.4 3.29 1.215 2.4 1.215 2.4 1 1.67 1 1.67 0.94 1.73 0.94 1.73 0.62 1.245 0.62 1.245 0.715 1.185 0.715 1.185 0.56 1.67 0.56 1.67 0.465 1.79 0.465 1.79 0.94 2.46 0.94 2.46 1.155 3.35 1.155 3.35 1.34 3.93 1.34 3.93 0.72 3.99 0.72 3.99 1.34 4.245 1.34 ;
      POLYGON 3.915 0.62 3.83 0.62 3.83 1.24 3.77 1.24 3.77 1.18 3.45 1.18 3.45 1.055 2.56 1.055 2.56 0.995 2.62 0.995 2.62 0.84 2.07 0.84 2.07 0.335 1.715 0.335 1.715 0.34 1.215 0.34 1.215 0.28 1.655 0.28 1.655 0.275 2.45 0.275 2.45 0.44 2.575 0.44 2.575 0.5 2.39 0.5 2.39 0.335 2.13 0.335 2.13 0.78 2.68 0.78 2.68 0.995 3.51 0.995 3.51 1.12 3.77 1.12 3.77 0.56 3.855 0.56 3.855 0.5 3.915 0.5 ;
      POLYGON 2.97 1.48 2.24 1.48 2.24 1.16 1.51 1.16 1.51 0.875 1.025 0.875 1.025 0.335 0.765 0.335 0.765 0.725 0.705 0.725 0.705 0.53 0.16 0.53 0.16 1.23 0.275 1.23 0.275 1.35 0.215 1.35 0.215 1.29 0.1 1.29 0.1 0.47 0.205 0.47 0.205 0.41 0.265 0.41 0.265 0.47 0.705 0.47 0.705 0.275 1.085 0.275 1.085 0.815 1.51 0.815 1.51 0.72 1.62 0.72 1.62 0.84 1.57 0.84 1.57 1.1 2.3 1.1 2.3 1.42 2.97 1.42 ;
      POLYGON 2.885 0.53 2.735 0.53 2.735 0.66 2.23 0.66 2.23 0.435 2.29 0.435 2.29 0.6 2.675 0.6 2.675 0.47 2.825 0.47 2.825 0.41 2.885 0.41 ;
      POLYGON 2.14 1.32 1.12 1.32 1.12 1.195 0.865 1.195 0.865 0.435 0.925 0.435 0.925 1.135 1.18 1.135 1.18 1.26 2.14 1.26 ;
  END
END DFFSRX4

MACRO DFFSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSRXL 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.47455 LAYER Metal1 ;
    ANTENNADIFFAREA 3.4816 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2268 LAYER Metal1 ;
      ANTENNAMAXAREACAR 15.31988525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 117.32804225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.635 0.945 0.635 0.945 1.315 0.885 1.315 0.885 0.73 0.86 0.73 0.86 0.6 0.885 0.6 0.885 0.575 0.94 0.575 0.94 0.515 1 0.515 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5291 LAYER Metal1 ;
    ANTENNADIFFAREA 3.4816 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2268 LAYER Metal1 ;
      ANTENNAMAXAREACAR 15.56040575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 118.5714285 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.315 1.02 0.235 1.02 0.235 0.73 0.06 0.73 0.06 0.6 0.235 0.6 0.235 0.54 0.315 0.54 ;
    END
  END QN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.26 0.755 6.34 1.255 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 0.925 5.66 0.925 5.66 0.485 5.74 0.485 5.74 0.79 5.8 0.79 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 32.68518525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.605 0.86 3.745 0.86 3.745 0.36 3.165 0.36 3.165 0.765 2.04 0.765 2.04 0.705 3.035 0.705 3.035 0.625 3.105 0.625 3.105 0.3 3.805 0.3 3.805 0.8 4.605 0.8 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 1.16 1.045 1.16 1.045 1.005 1.195 1.005 1.195 0.9 1.365 0.9 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 1.77 0 1.77 0 1.65 0.49 1.65 0.49 1.01 0.55 1.01 0.55 1.65 1.15 1.65 1.15 1.29 1.21 1.29 1.21 1.65 1.86 1.65 1.86 1.54 1.98 1.54 1.98 1.65 2.56 1.65 2.56 1.205 2.62 1.205 2.62 1.65 4.105 1.65 4.105 1.54 4.225 1.54 4.225 1.65 4.705 1.65 4.705 1.54 4.825 1.54 4.825 1.65 5.735 1.65 5.735 1.51 5.795 1.51 5.795 1.65 6.44 1.65 6.44 1.02 6.5 1.02 6.5 1.65 6.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 0.06 6.395 0.06 6.395 0.635 6.335 0.635 6.335 0.06 5.755 0.06 5.755 0.385 5.695 0.385 5.695 0.06 4.825 0.06 4.825 0.17 4.705 0.17 4.705 0.06 1.99 0.06 1.99 0.445 1.93 0.445 1.93 0.06 1.205 0.06 1.205 0.635 1.145 0.635 1.145 0.06 0.52 0.06 0.52 0.635 0.46 0.635 0.46 0.06 0 0.06 0 -0.06 6.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.16 1.305 5.635 1.305 5.635 1.34 3.325 1.34 3.325 1.28 5.575 1.28 5.575 1.245 6.1 1.245 6.1 0.54 6.16 0.54 ;
      POLYGON 5.96 1.145 5.9 1.145 5.9 1.085 5.475 1.085 5.475 1.18 3.225 1.18 3.225 1.265 3.085 1.265 3.085 1.205 3.165 1.205 3.165 1.12 3.425 1.12 3.425 0.74 3.485 0.74 3.485 1.12 5.035 1.12 5.035 0.63 5.095 0.63 5.095 1.12 5.415 1.12 5.415 0.74 5.475 0.74 5.475 1.025 5.9 1.025 5.9 0.29 5.96 0.29 ;
      POLYGON 5.315 1.02 5.195 1.02 5.195 0.35 4.43 0.35 4.43 0.29 5.255 0.29 5.255 0.96 5.315 0.96 ;
      POLYGON 4.925 0.765 4.865 0.765 4.865 0.7 4.765 0.7 4.765 1.02 3.585 1.02 3.585 0.46 3.645 0.46 3.645 0.96 4.705 0.96 4.705 0.7 4.11 0.7 4.11 0.475 4.17 0.475 4.17 0.64 4.925 0.64 ;
      POLYGON 4.565 0.54 4.27 0.54 4.27 0.375 3.965 0.375 3.965 0.57 3.905 0.57 3.905 0.315 4.33 0.315 4.33 0.48 4.565 0.48 ;
      POLYGON 3.44 0.64 3.325 0.64 3.325 0.925 3.24 0.925 3.24 1.02 3.18 1.02 3.18 0.925 1.88 0.925 1.88 0.715 1.94 0.715 1.94 0.865 3.265 0.865 3.265 0.58 3.38 0.58 3.38 0.46 3.44 0.46 ;
      RECT 2.095 1.025 3.065 1.105 ;
      POLYGON 3.005 0.525 2.935 0.525 2.935 0.595 2.455 0.595 2.455 0.445 2.415 0.445 2.415 0.365 2.535 0.365 2.535 0.515 2.855 0.515 2.855 0.445 3.005 0.445 ;
      POLYGON 2.755 0.415 2.635 0.415 2.635 0.265 2.28 0.265 2.28 0.445 2.2 0.445 2.2 0.185 2.715 0.185 2.715 0.335 2.755 0.335 ;
      POLYGON 2.46 1.265 1.525 1.265 1.525 1.325 1.465 1.325 1.465 0.54 1.525 0.54 1.525 1.205 2.46 1.205 ;
      POLYGON 2.355 0.605 1.78 0.605 1.78 1.02 1.72 1.02 1.72 0.41 1.365 0.41 1.365 0.8 1.045 0.8 1.045 0.74 1.305 0.74 1.305 0.35 1.78 0.35 1.78 0.545 2.355 0.545 ;
      POLYGON 0.785 1.02 0.705 1.02 0.705 0.91 0.67 0.91 0.67 0.815 0.415 0.815 0.415 0.735 0.67 0.735 0.67 0.54 0.75 0.54 0.75 0.83 0.785 0.83 ;
  END
END DFFSRXL

MACRO DFFSX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSX1 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6114 LAYER Metal1 ;
    ANTENNADIFFAREA 2.622225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2205 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.843084 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 91.6190475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.65 0.36 0.73 1.29 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6114 LAYER Metal1 ;
    ANTENNADIFFAREA 2.622225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2205 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.843084 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 91.6190475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.05 0.42 0.13 1.29 ;
    END
  END QN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.9814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.07 0.555 4.15 0.96 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.35185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.87 0.555 3.95 0.98 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.074074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.765 0.99 1.52 0.99 1.52 0.895 1.5 0.895 1.5 0.815 1.765 0.815 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.305 1.65 0.305 1.285 0.365 1.285 0.365 1.65 0.875 1.65 0.875 0.995 0.935 0.995 0.935 1.65 1.25 1.65 1.25 1.09 1.31 1.09 1.31 1.65 1.69 1.65 1.69 1.465 1.81 1.465 1.81 1.65 2.1 1.65 2.1 1.465 2.22 1.465 2.22 1.65 3.175 1.65 3.175 1.465 3.3 1.465 3.3 1.65 3.96 1.65 3.96 1.08 4.02 1.08 4.02 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 4.11 0.06 4.11 0.24 4.05 0.24 4.05 0.06 3.29 0.06 3.29 0.26 3.17 0.26 3.17 0.06 1.785 0.06 1.785 0.2 1.725 0.2 1.725 0.06 0.97 0.06 0.97 0.28 0.91 0.28 0.91 0.06 0.365 0.06 0.365 0.33 0.305 0.33 0.305 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.28 1.12 4.225 1.12 4.225 1.18 4.165 1.18 4.165 1.06 4.22 1.06 4.22 0.415 3.61 0.415 3.61 0.935 3.55 0.935 3.55 0.415 2.69 0.415 2.69 0.925 2.63 0.925 2.63 0.415 2.385 0.415 2.385 0.355 4.28 0.355 ;
      POLYGON 3.77 1.095 3.685 1.095 3.685 1.405 1.94 1.405 1.94 1.345 3.625 1.345 3.625 1.035 3.71 1.035 3.71 0.515 3.77 0.515 ;
      POLYGON 3.45 0.935 3.39 0.935 3.39 0.755 2.985 0.755 2.985 1.015 3.045 1.015 3.045 1.075 2.925 1.075 2.925 0.49 3.01 0.49 3.01 0.695 3.45 0.695 ;
      POLYGON 3.29 0.915 3.205 0.915 3.205 1.245 2.38 1.245 2.38 0.98 2.075 0.98 2.075 1.085 1.865 1.085 1.865 1.025 1.98 1.025 1.98 0.515 2.075 0.515 2.075 0.92 2.44 0.92 2.44 1.185 2.705 1.185 2.705 1.025 2.75 1.025 2.75 0.515 2.81 0.515 2.81 1.085 2.765 1.085 2.765 1.185 3.145 1.185 3.145 0.855 3.29 0.855 ;
      POLYGON 2.56 1.095 2.5 1.095 2.5 0.785 2.135 0.785 2.135 0.44 1.57 0.44 1.57 0.745 1.035 0.745 1.035 0.685 1.51 0.685 1.51 0.38 2.195 0.38 2.195 0.725 2.495 0.725 2.495 0.605 2.435 0.605 2.435 0.545 2.56 0.545 ;
      POLYGON 2.32 0.625 2.26 0.625 2.26 0.32 1.37 0.32 1.37 0.58 1.25 0.58 1.25 0.52 1.31 0.52 1.31 0.26 2.32 0.26 ;
      POLYGON 2.32 1.245 1.485 1.245 1.485 1.09 1.545 1.09 1.545 1.185 2.26 1.185 2.26 1.06 2.32 1.06 ;
      POLYGON 1.42 0.925 1.36 0.925 1.36 0.935 1.14 0.935 1.14 1.02 1.08 1.02 1.08 0.935 0.91 0.935 0.91 0.74 0.79 0.74 0.79 0.68 0.91 0.68 0.91 0.495 1.17 0.495 1.17 0.555 0.97 0.555 0.97 0.875 1.3 0.875 1.3 0.865 1.42 0.865 ;
      POLYGON 0.53 1.02 0.45 1.02 0.45 0.81 0.195 0.81 0.195 0.73 0.45 0.73 0.45 0.54 0.53 0.54 ;
  END
END DFFSX1

MACRO DFFSX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSX2 0 0 ;
  SIZE 6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3152 LAYER Metal1 ;
    ANTENNADIFFAREA 3.57945 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.285975 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.59262175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 90.59533175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.35 0.65 5.34 0.65 5.34 1.29 5.26 1.29 5.26 0.65 5.23 0.65 5.23 0.57 5.35 0.57 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3152 LAYER Metal1 ;
    ANTENNADIFFAREA 3.57945 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.285975 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.59262175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 90.59533175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.74 1.29 4.66 1.29 4.66 0.63 4.62 0.63 4.62 0.55 4.74 0.55 ;
    END
  END Q
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.46 0.75 3.54 1.25 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.61 0.34 1.11 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 1.77 0 1.77 0 1.65 0.41 1.65 0.41 1.21 0.47 1.21 0.47 1.65 1.13 1.65 1.13 1.51 1.19 1.51 1.19 1.65 2.91 1.65 2.91 1.54 3.03 1.54 3.03 1.65 3.435 1.65 3.435 1.51 3.495 1.51 3.495 1.65 3.805 1.65 3.805 1.51 3.865 1.51 3.865 1.65 4.45 1.65 4.45 1.12 4.51 1.12 4.51 1.65 4.905 1.65 4.905 0.92 4.965 0.92 4.965 1.65 5.465 1.65 5.465 0.995 5.525 0.995 5.525 1.65 6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 0.06 5.585 0.06 5.585 0.17 5.465 0.17 5.465 0.06 5.025 0.06 5.025 0.17 4.905 0.17 4.905 0.06 4.505 0.06 4.505 0.17 4.385 0.17 4.385 0.06 3.455 0.06 3.455 0.33 3.335 0.33 3.335 0.27 3.395 0.27 3.395 0.06 1.495 0.06 1.495 0.17 1.375 0.17 1.375 0.06 0.5 0.06 0.5 0.2 0.44 0.2 0.44 0.06 0 0.06 0 -0.06 6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.805 0.63 5.775 0.63 5.775 1.02 5.715 1.02 5.715 0.81 5.44 0.81 5.44 0.75 5.715 0.75 5.715 0.63 5.685 0.63 5.685 0.57 5.805 0.57 ;
      POLYGON 5.745 0.45 4.9 0.45 4.9 0.82 4.84 0.82 4.84 0.45 4.5 0.45 4.5 0.73 4.56 0.73 4.56 0.79 4.5 0.79 4.5 1.02 4.335 1.02 4.335 1.07 4.215 1.07 4.215 1.01 4.275 1.01 4.275 0.96 4.44 0.96 4.44 0.7 3.8 0.7 3.8 0.64 4.18 0.64 4.18 0.54 4.24 0.54 4.24 0.64 4.44 0.64 4.44 0.39 5.685 0.39 5.685 0.33 5.745 0.33 ;
      POLYGON 4.335 0.86 3.64 0.86 3.64 0.65 3.195 0.65 3.195 0.83 2.9 0.83 2.9 0.77 3.135 0.77 3.135 0.59 3.7 0.59 3.7 0.8 4.335 0.8 ;
      POLYGON 3.935 0.49 3.16 0.49 3.16 0.355 2.64 0.355 2.64 0.57 2.335 0.57 2.335 0.51 2.58 0.51 2.58 0.295 3.22 0.295 3.22 0.43 3.935 0.43 ;
      POLYGON 3.7 1.41 3.3 1.41 3.3 1.265 3.015 1.265 3.015 1.205 2.48 1.205 2.48 1.145 3.075 1.145 3.075 1.205 3.36 1.205 3.36 1.35 3.64 1.35 3.64 1.03 3.7 1.03 ;
      POLYGON 3.235 1.105 3.175 1.105 3.175 1.045 2.38 1.045 2.38 1.365 1.45 1.365 1.45 1.01 1.34 1.01 1.34 0.95 1.51 0.95 1.51 1.305 1.925 1.305 1.925 1.175 1.84 1.175 1.84 0.505 1.9 0.505 1.9 1.115 1.985 1.115 1.985 1.305 2.32 1.305 2.32 0.985 2.74 0.985 2.74 0.455 3.06 0.455 3.06 0.515 2.8 0.515 2.8 0.985 3.235 0.985 ;
      POLYGON 3.2 1.425 2.54 1.425 2.54 1.525 1.29 1.525 1.29 1.235 0.945 1.235 0.945 1.175 0.86 1.175 0.86 0.505 0.8 0.505 0.8 0.445 0.92 0.445 0.92 1.115 1.005 1.115 1.005 1.175 1.35 1.175 1.35 1.465 2.48 1.465 2.48 1.365 3.2 1.365 ;
      POLYGON 2.58 0.885 2.22 0.885 2.22 1.11 2.1 1.11 2.1 1.05 2.16 1.05 2.16 0.505 2.22 0.505 2.22 0.825 2.58 0.825 ;
      POLYGON 2.325 0.22 2.06 0.22 2.06 0.915 2 0.915 2 0.31 1.51 0.31 1.51 0.345 1.08 0.345 1.08 0.955 1.02 0.955 1.02 0.345 0.7 0.345 0.7 0.725 0.64 0.725 0.64 0.51 0.16 0.51 0.16 1.21 0.265 1.21 0.265 1.33 0.205 1.33 0.205 1.27 0.1 1.27 0.1 0.45 0.205 0.45 0.205 0.39 0.265 0.39 0.265 0.45 0.64 0.45 0.64 0.285 1.45 0.285 1.45 0.25 2 0.25 2 0.16 2.325 0.16 ;
      POLYGON 1.74 0.81 1.73 0.81 1.73 1.205 1.61 1.205 1.61 1.145 1.67 1.145 1.67 0.75 1.18 0.75 1.18 0.69 1.61 0.69 1.61 0.445 1.73 0.445 1.73 0.505 1.67 0.505 1.67 0.69 1.74 0.69 ;
  END
END DFFSX2

MACRO DFFSX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSX4 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4585 LAYER Metal1 ;
    ANTENNADIFFAREA 4.0829 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4392 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.87454475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 60.976776 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.79 0.66 5.34 0.66 5.34 0.94 5.73 0.94 5.73 1.33 5.67 1.33 5.67 1 5.32 1 5.32 1.33 5.26 1.33 5.26 0.54 5.32 0.54 5.32 0.6 5.73 0.6 5.73 0.54 5.79 0.54 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4585 LAYER Metal1 ;
    ANTENNADIFFAREA 4.0829 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4392 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.87454475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 60.976776 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.91 1.33 4.85 1.33 4.85 1 4.5 1 4.5 1.33 4.44 1.33 4.44 0.94 4.46 0.94 4.46 0.625 4.32 0.625 4.32 0.505 4.38 0.505 4.38 0.565 4.79 0.565 4.79 0.505 4.85 0.505 4.85 0.625 4.52 0.625 4.52 0.79 4.54 0.79 4.54 0.94 4.91 0.94 ;
    END
  END Q
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 22.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.575 0.97 3.515 0.97 3.515 0.91 3.14 0.91 3.14 0.92 3.06 0.92 3.06 0.79 3.08 0.79 3.08 0.395 2.32 0.395 2.32 0.44 1.94 0.44 1.94 0.435 1.82 0.435 1.82 0.375 2 0.375 2 0.38 2.26 0.38 2.26 0.335 3.14 0.335 3.14 0.85 3.575 0.85 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.655 0.895 0.54 0.895 0.54 0.995 0.46 0.995 0.46 0.775 0.575 0.775 0.575 0.61 0.655 0.61 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.36 1.09 0.28 1.09 0.28 0.96 0.26 0.96 0.26 0.61 0.36 0.61 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 1.77 0 1.77 0 1.65 0.505 1.65 0.505 1.095 0.565 1.095 0.565 1.65 1.335 1.65 1.335 1.51 1.395 1.51 1.395 1.65 1.825 1.65 1.825 1.54 1.945 1.54 1.945 1.65 3.22 1.65 3.22 1.49 3.34 1.49 3.34 1.55 3.28 1.55 3.28 1.65 3.675 1.65 3.675 1.24 3.795 1.24 3.795 1.3 3.735 1.3 3.735 1.65 4.235 1.65 4.235 0.945 4.295 0.945 4.295 1.65 4.645 1.65 4.645 1.1 4.705 1.1 4.705 1.65 5.055 1.65 5.055 0.94 5.115 0.94 5.115 1.65 5.465 1.65 5.465 1.1 5.525 1.1 5.525 1.65 5.875 1.65 5.875 1.1 5.935 1.1 5.935 1.65 6.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 0.06 6.11 0.06 6.11 0.52 6.05 0.52 6.05 0.06 5.585 0.06 5.585 0.17 5.465 0.17 5.465 0.06 5.115 0.06 5.115 0.17 4.995 0.17 4.995 0.06 4.645 0.06 4.645 0.17 4.525 0.17 4.525 0.06 4.06 0.06 4.06 0.575 4 0.575 4 0.06 3.65 0.06 3.65 0.59 3.59 0.59 3.59 0.06 2.16 0.06 2.16 0.28 2.1 0.28 2.1 0.06 1.46 0.06 1.46 0.17 1.34 0.17 1.34 0.06 0.5 0.06 0.5 0.35 0.44 0.35 0.44 0.06 0 0.06 0 -0.06 6.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.315 1 6.14 1 6.14 1.33 6.08 1.33 6.08 1 5.83 1 5.83 0.78 5.89 0.78 5.89 0.94 6.255 0.94 6.255 0.54 6.315 0.54 ;
      POLYGON 6.075 0.84 6.015 0.84 6.015 0.68 5.89 0.68 5.89 0.405 4.22 0.405 4.22 0.725 4.36 0.725 4.36 0.845 4.3 0.845 4.3 0.785 4.06 0.785 4.06 1.33 4 1.33 4 0.75 3.315 0.75 3.315 0.69 3.795 0.69 3.795 0.54 3.855 0.54 3.855 0.69 4.16 0.69 4.16 0.345 5.95 0.345 5.95 0.62 6.075 0.62 ;
      POLYGON 3.9 0.97 3.735 0.97 3.735 1.13 2.68 1.13 2.68 1.225 2.62 1.225 2.62 1.07 2.9 1.07 2.9 0.495 2.96 0.495 2.96 1.07 3.675 1.07 3.675 0.91 3.84 0.91 3.84 0.85 3.9 0.85 ;
      RECT 2.795 1.23 3.575 1.31 ;
      POLYGON 2.8 0.97 2.47 0.97 2.47 1.31 2.41 1.31 2.41 1.25 1.9 1.25 1.9 1.145 1.62 1.145 1.62 0.755 1.235 0.755 1.235 0.695 1.5 0.695 1.5 0.53 1.56 0.53 1.56 0.695 1.68 0.695 1.68 1.085 1.96 1.085 1.96 1.19 2.41 1.19 2.41 0.91 2.74 0.91 2.74 0.585 2.665 0.585 2.665 0.525 2.8 0.525 ;
      POLYGON 2.64 0.81 2.18 0.81 2.18 1.09 2.06 1.09 2.06 1.03 2.12 1.03 2.12 0.81 1.78 0.81 1.78 0.595 1.66 0.595 1.66 0.43 1.135 0.43 1.135 0.545 1.075 0.545 1.075 0.37 1.72 0.37 1.72 0.535 1.84 0.535 1.84 0.75 2.42 0.75 2.42 0.53 2.48 0.53 2.48 0.75 2.58 0.75 2.58 0.69 2.64 0.69 ;
      POLYGON 2.105 1.41 1.05 1.41 1.05 1.495 0.99 1.495 0.99 1.41 0.755 1.41 0.755 0.51 0.135 0.51 0.135 1.215 0.075 1.215 0.075 0.45 0.235 0.45 0.235 0.255 0.295 0.255 0.295 0.45 0.815 0.45 0.815 1.35 2.105 1.35 ;
      POLYGON 1.52 0.925 0.975 0.925 0.975 1.12 0.915 1.12 0.915 0.255 0.975 0.255 0.975 0.865 1.52 0.865 ;
  END
END DFFSX4

MACRO DFFSXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFSXL 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.696275 LAYER Metal1 ;
    ANTENNADIFFAREA 2.785575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1944 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.86972725 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 107.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.49 0.94 1.02 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.696275 LAYER Metal1 ;
    ANTENNADIFFAREA 2.785575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1944 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.86972725 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 107.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.305 1.02 0.225 1.02 0.225 0.73 0.06 0.73 0.06 0.6 0.225 0.6 0.225 0.54 0.305 0.54 ;
    END
  END QN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.66 0.46 4.74 0.96 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.46 0.46 4.54 0.96 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.185 0.94 2.035 0.94 2.035 0.895 1.73 0.895 1.73 0.815 2.185 0.815 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 1.77 0 1.77 0 1.65 0.515 1.65 0.515 1.285 0.575 1.285 0.575 1.65 1.15 1.65 1.15 1.285 1.21 1.285 1.21 1.65 1.515 1.65 1.515 1.06 1.575 1.06 1.575 1.65 2.08 1.65 2.08 1.295 2.14 1.295 2.14 1.65 2.52 1.65 2.52 1.54 2.64 1.54 2.64 1.65 4.055 1.65 4.055 1.51 4.115 1.51 4.115 1.65 4.55 1.65 4.55 1.06 4.61 1.06 4.61 1.65 5 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 0.06 4.7 0.06 4.7 0.2 4.64 0.2 4.64 0.06 3.88 0.06 3.88 0.17 3.76 0.17 3.76 0.06 1.945 0.06 1.945 0.2 1.885 0.2 1.885 0.06 1.21 0.06 1.21 0.2 1.15 0.2 1.15 0.06 0.575 0.06 0.575 0.2 0.515 0.2 0.515 0.06 0 0.06 0 -0.06 5 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.9 1.12 4.815 1.12 4.815 1.18 4.755 1.18 4.755 1.06 4.84 1.06 4.84 0.36 4.2 0.36 4.2 0.915 4.14 0.915 4.14 0.385 3.255 0.385 3.255 0.895 3.195 0.895 3.195 0.385 3.165 0.385 3.165 0.38 3.08 0.38 3.08 0.32 3.2 0.32 3.2 0.325 4.14 0.325 4.14 0.3 4.335 0.3 4.335 0.16 4.455 0.16 4.455 0.3 4.9 0.3 ;
      POLYGON 4.36 1.075 4.275 1.075 4.275 1.135 3.955 1.135 3.955 1.375 2.36 1.375 2.36 1.315 3.895 1.315 3.895 1.075 4.215 1.075 4.215 1.015 4.3 1.015 4.3 0.495 4.36 0.495 ;
      POLYGON 4.04 0.915 3.98 0.915 3.98 0.735 3.575 0.735 3.575 0.995 3.635 0.995 3.635 1.055 3.515 1.055 3.515 0.68 3.525 0.68 3.525 0.515 3.645 0.515 3.645 0.575 3.585 0.575 3.585 0.675 4.04 0.675 ;
      POLYGON 3.88 0.895 3.795 0.895 3.795 1.215 2.875 1.215 2.875 0.96 2.405 0.96 2.405 1.035 2.285 1.035 2.285 0.975 2.345 0.975 2.345 0.9 2.44 0.9 2.44 0.49 2.5 0.49 2.5 0.9 2.935 0.9 2.935 1.155 3.27 1.155 3.27 0.995 3.355 0.995 3.355 0.485 3.415 0.485 3.415 1.055 3.33 1.055 3.33 1.155 3.735 1.155 3.735 0.835 3.88 0.835 ;
      POLYGON 3.155 1.055 3.035 1.055 3.035 0.785 2.6 0.785 2.6 0.39 2.34 0.39 2.34 0.48 2.265 0.48 2.265 0.715 1.32 0.715 1.32 0.775 1.26 0.775 1.26 0.655 2.205 0.655 2.205 0.42 2.28 0.42 2.28 0.33 2.66 0.33 2.66 0.725 3.035 0.725 3.035 0.575 2.975 0.575 2.975 0.515 3.095 0.515 3.095 0.995 3.155 0.995 ;
      POLYGON 2.875 0.625 2.795 0.625 2.795 0.35 2.76 0.35 2.76 0.16 2.84 0.16 2.84 0.27 2.875 0.27 ;
      POLYGON 2.775 1.12 2.565 1.12 2.565 1.195 1.845 1.195 1.845 1.04 1.905 1.04 1.905 1.135 2.505 1.135 2.505 1.06 2.775 1.06 ;
      POLYGON 2.18 0.32 2.105 0.32 2.105 0.555 1.515 0.555 1.515 0.495 2.045 0.495 2.045 0.26 2.18 0.26 ;
      POLYGON 1.63 0.875 1.48 0.875 1.48 0.935 1.375 0.935 1.375 1.02 1.315 1.02 1.315 0.935 1.1 0.935 1.1 0.74 1.04 0.74 1.04 0.68 1.1 0.68 1.1 0.495 1.405 0.495 1.405 0.555 1.16 0.555 1.16 0.875 1.42 0.875 1.42 0.815 1.63 0.815 ;
      POLYGON 0.74 1.02 0.66 1.02 0.66 0.81 0.405 0.81 0.405 0.73 0.66 0.73 0.66 0.54 0.74 0.54 ;
  END
END DFFSXL

MACRO DFFTRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFTRX1 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.54155 LAYER Metal1 ;
    ANTENNADIFFAREA 2.729575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2205 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.52630375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 88.462585 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.975 0.53 0.94 0.53 0.94 0.89 0.96 0.89 0.96 1.34 0.9 1.34 0.9 0.95 0.88 0.95 0.88 0.54 0.86 0.54 0.86 0.41 0.975 0.41 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.54155 LAYER Metal1 ;
    ANTENNADIFFAREA 2.729575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2205 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.52630375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 88.462585 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.325 1.29 0.245 1.29 0.245 0.73 0.06 0.73 0.06 0.6 0.245 0.6 0.245 0.54 0.325 0.54 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.46 0.365 4.54 0.865 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.32 1.005 4.24 1.005 4.24 0.87 4.14 0.87 4.14 0.92 4.06 0.92 4.06 0.79 4.24 0.79 4.24 0.735 4.32 0.735 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.29629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 1.06 1.14 1.06 1.14 1.11 1.06 1.11 1.06 0.98 1.26 0.98 1.26 0.78 1.34 0.78 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.47 1.65 0.47 0.995 0.53 0.995 0.53 1.65 1.105 1.65 1.105 1.22 1.165 1.22 1.165 1.65 2.03 1.65 2.03 1.49 2.15 1.49 2.15 1.55 2.09 1.55 2.09 1.65 3.02 1.65 3.02 1.49 3.14 1.49 3.14 1.55 3.08 1.55 3.08 1.65 4.105 1.65 4.105 1.51 4.165 1.51 4.165 1.65 4.625 1.65 4.625 1.125 4.685 1.125 4.685 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 4.205 0.06 4.205 0.635 4.145 0.635 4.145 0.06 3.14 0.06 3.14 0.17 3.02 0.17 3.02 0.06 2.09 0.06 2.09 0.61 2.03 0.61 2.03 0.06 1.18 0.06 1.18 0.52 1.12 0.52 1.12 0.06 0.56 0.06 0.56 0.2 0.5 0.2 0.5 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.7 1.025 4.48 1.025 4.48 1.375 3.615 1.375 3.615 0.995 3.74 0.995 3.74 0.515 3.8 0.515 3.8 1.055 3.675 1.055 3.675 1.315 4.42 1.315 4.42 0.965 4.64 0.965 4.64 0.54 4.7 0.54 ;
      POLYGON 4 0.69 3.96 0.69 3.96 1.215 3.84 1.215 3.84 1.155 3.9 1.155 3.9 0.63 3.94 0.63 3.94 0.53 3.9 0.53 3.9 0.415 3.64 0.415 3.64 0.895 3.52 0.895 3.52 0.835 3.58 0.835 3.58 0.415 2.685 0.415 2.685 0.705 2.745 0.705 2.745 0.825 2.685 0.825 2.685 0.875 2.48 0.875 2.48 0.935 2.42 0.935 2.42 0.815 2.625 0.815 2.625 0.355 3.285 0.355 3.285 0.275 3.405 0.275 3.405 0.355 3.96 0.355 3.96 0.47 4 0.47 ;
      POLYGON 3.48 0.605 3.42 0.605 3.42 0.995 3.47 0.995 3.47 1.16 3.41 1.16 3.41 1.055 3.36 1.055 3.36 0.925 3.005 0.925 3.005 0.865 3.36 0.865 3.36 0.545 3.48 0.545 ;
      POLYGON 3.435 1.385 1.44 1.385 1.44 0.54 1.5 0.54 1.5 1.325 3.435 1.325 ;
      POLYGON 3.235 0.765 2.905 0.765 2.905 1.13 2.785 1.13 2.785 1.07 2.845 1.07 2.845 0.605 2.785 0.605 2.785 0.545 2.905 0.545 2.905 0.705 3.235 0.705 ;
      POLYGON 2.585 1.13 2.26 1.13 2.26 0.93 1.96 0.93 1.96 0.99 1.9 0.99 1.9 0.87 2.26 0.87 2.26 0.655 2.465 0.655 2.465 0.515 2.525 0.515 2.525 0.715 2.32 0.715 2.32 1.07 2.585 1.07 ;
      POLYGON 2.16 0.77 1.8 0.77 1.8 1.09 1.915 1.09 1.915 1.15 1.74 1.15 1.74 0.55 1.825 0.55 1.825 0.45 1.6 0.45 1.6 0.44 1.34 0.44 1.34 0.68 1.16 0.68 1.16 0.79 1.04 0.79 1.04 0.62 1.28 0.62 1.28 0.38 1.66 0.38 1.66 0.39 1.885 0.39 1.885 0.61 1.8 0.61 1.8 0.71 2.16 0.71 ;
      POLYGON 0.76 1.02 0.68 1.02 0.68 0.85 0.425 0.85 0.425 0.77 0.68 0.77 0.68 0.54 0.76 0.54 ;
  END
END DFFTRX1

MACRO DFFTRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFTRX2 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.652525 LAYER Metal1 ;
    ANTENNADIFFAREA 2.959675 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.285975 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.27537375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 72.027275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.25 0.65 4.17 0.65 4.17 0.88 4.19 0.88 4.19 1.29 4.11 1.29 4.11 0.94 4.09 0.94 4.09 0.73 4.06 0.73 4.06 0.6 4.09 0.6 4.09 0.57 4.25 0.57 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.652525 LAYER Metal1 ;
    ANTENNADIFFAREA 2.959675 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.285975 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.27537375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 72.027275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.78 1.29 3.72 1.29 3.72 0.73 3.66 0.73 3.66 0.57 3.78 0.57 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 0.895 3.18 0.895 3.18 0.77 3.26 0.77 3.26 0.535 3.34 0.535 3.34 0.77 3.4 0.77 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.2 1.015 0.12 1.015 0.12 0.73 0.06 0.73 0.06 0.575 0.2 0.575 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.095 1.65 0.095 1.115 0.155 1.115 0.155 1.65 0.54 1.65 0.54 1.405 0.6 1.405 0.6 1.65 1.58 1.65 1.58 1.54 1.7 1.54 1.7 1.65 2.63 1.65 2.63 1.49 2.75 1.49 2.75 1.55 2.69 1.55 2.69 1.65 3.515 1.65 3.515 0.92 3.575 0.92 3.575 1.65 3.925 1.65 3.925 0.945 3.985 0.945 3.985 1.65 4.335 1.65 4.335 0.91 4.395 0.91 4.395 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 4.455 0.06 4.455 0.2 4.395 0.2 4.395 0.06 4.015 0.06 4.015 0.17 3.895 0.17 3.895 0.06 3.545 0.06 3.545 0.17 3.425 0.17 3.425 0.06 2.68 0.06 2.68 0.575 2.62 0.575 2.62 0.06 1.64 0.06 1.64 0.16 1.7 0.16 1.7 0.22 1.58 0.22 1.58 0.06 0.535 0.06 0.535 0.475 0.475 0.475 0.475 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.69 0.81 4.63 0.81 4.63 1.02 4.57 1.02 4.57 0.81 4.27 0.81 4.27 0.75 4.63 0.75 4.63 0.54 4.69 0.54 ;
      POLYGON 4.675 0.435 3.94 0.435 3.94 0.845 3.88 0.845 3.88 0.435 3.56 0.435 3.56 0.82 3.5 0.82 3.5 0.435 2.885 0.435 2.885 0.58 2.92 0.58 2.92 1.155 2.985 1.155 2.985 1.215 2.86 1.215 2.86 1.01 2.66 1.01 2.66 0.89 2.72 0.89 2.72 0.95 2.86 0.95 2.86 0.645 2.825 0.645 2.825 0.375 4.675 0.375 ;
      POLYGON 3.305 1.39 2.475 1.39 2.475 1.405 1.295 1.405 1.295 1.345 2.43 1.345 2.43 1.33 3.245 1.33 3.245 1.055 3.02 1.055 3.02 0.57 3.16 0.57 3.16 0.63 3.08 0.63 3.08 0.995 3.305 0.995 ;
      POLYGON 2.76 0.79 2.56 0.79 2.56 1.12 2.33 1.12 2.33 1.18 2.27 1.18 2.27 1.06 2.5 1.06 2.5 0.79 2.28 0.79 2.28 0.54 2.34 0.54 2.34 0.73 2.76 0.73 ;
      POLYGON 2.4 0.95 2.12 0.95 2.12 0.88 2.035 0.88 2.035 0.76 2.12 0.76 2.12 0.44 1.1 0.44 1.1 0.87 1.16 0.87 1.16 0.93 1.04 0.93 1.04 0.44 0.74 0.44 0.74 0.54 0.765 0.54 0.765 1.14 0.705 1.14 0.705 0.6 0.68 0.6 0.68 0.38 1.3 0.38 1.3 0.305 1.42 0.305 1.42 0.38 2.18 0.38 2.18 0.89 2.4 0.89 ;
      POLYGON 2.02 0.66 1.935 0.66 1.935 1.18 1.875 1.18 1.875 0.99 1.485 0.99 1.485 0.93 1.875 0.93 1.875 0.6 1.96 0.6 1.96 0.54 2.02 0.54 ;
      POLYGON 1.775 0.8 1.32 0.8 1.32 1.18 1.26 1.18 1.26 0.63 1.2 0.63 1.2 0.57 1.32 0.57 1.32 0.74 1.775 0.74 ;
      POLYGON 1.115 1.3 0.3 1.3 0.3 0.475 0.165 0.475 0.165 0.355 0.225 0.355 0.225 0.415 0.36 0.415 0.36 1.24 0.88 1.24 0.88 0.54 0.94 0.54 0.94 1.155 1.115 1.155 ;
  END
END DFFTRX2

MACRO DFFTRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFTRX4 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.40535 LAYER Metal1 ;
    ANTENNADIFFAREA 3.8476 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4392 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.75352925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 59.5286885 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.66 0.545 5.14 0.545 5.14 0.9 5.55 0.9 5.55 1.29 5.49 1.29 5.49 0.96 5.14 0.96 5.14 1.29 5.06 1.29 5.06 0.79 5.07 0.79 5.07 0.485 5.66 0.485 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.40535 LAYER Metal1 ;
    ANTENNADIFFAREA 3.8476 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4392 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.75352925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 59.5286885 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.73 1.29 4.67 1.29 4.67 0.96 4.32 0.96 4.32 1.29 4.26 1.29 4.26 0.79 4.28 0.79 4.28 0.545 4.13 0.545 4.13 0.485 4.72 0.485 4.72 0.545 4.34 0.545 4.34 0.9 4.73 0.9 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.435 0.895 1.125 0.895 1.125 0.625 1.42 0.625 1.42 0.815 1.435 0.815 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 1.055 0.325 1.055 0.325 0.69 0.405 0.69 0.405 0.79 0.54 0.79 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.225 1.055 0.14 1.055 0.14 1.11 0.06 1.11 0.06 0.98 0.095 0.98 0.095 0.695 0.225 0.695 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 1.77 0 1.77 0 1.65 0.13 1.65 0.13 1.51 0.19 1.51 0.19 1.65 0.53 1.65 0.53 1.315 0.59 1.315 0.59 1.65 1.53 1.65 1.53 1.315 1.59 1.315 1.59 1.65 2.545 1.65 2.545 1.075 2.605 1.075 2.605 1.65 3.615 1.65 3.615 1.03 3.675 1.03 3.675 1.65 4.055 1.65 4.055 0.97 4.115 0.97 4.115 1.65 4.465 1.65 4.465 1.06 4.525 1.06 4.525 1.65 4.875 1.65 4.875 0.9 4.935 0.9 4.935 1.65 5.285 1.65 5.285 1.06 5.345 1.06 5.345 1.65 5.72 1.65 5.72 1.02 5.78 1.02 5.78 1.65 6.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 0.06 5.98 0.06 5.98 0.435 5.92 0.435 5.92 0.06 5.425 0.06 5.425 0.17 5.305 0.17 5.305 0.06 4.955 0.06 4.955 0.17 4.835 0.17 4.835 0.06 4.485 0.06 4.485 0.17 4.365 0.17 4.365 0.06 4.015 0.06 4.015 0.17 3.895 0.17 3.895 0.06 3.545 0.06 3.545 0.55 3.485 0.55 3.485 0.06 2.665 0.06 2.665 0.17 2.545 0.17 2.545 0.06 1.485 0.06 1.485 0.365 1.425 0.365 1.425 0.06 0.175 0.06 0.175 0.59 0.115 0.59 0.115 0.06 0 0.06 0 -0.06 6.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.185 0.595 6.09 0.595 6.09 0.92 5.985 0.92 5.985 1.29 5.925 1.29 5.925 0.92 5.65 0.92 5.65 0.77 5.77 0.77 5.77 0.86 6.03 0.86 6.03 0.535 6.125 0.535 6.125 0.455 6.185 0.455 ;
      POLYGON 5.93 0.76 5.87 0.76 5.87 0.67 5.76 0.67 5.76 0.385 3.75 0.385 3.75 0.485 4.005 0.485 4.005 0.77 4.155 0.77 4.155 0.87 3.88 0.87 3.88 1.29 3.82 1.29 3.82 0.87 3.645 0.87 3.645 0.93 3.585 0.93 3.585 0.81 3.945 0.81 3.945 0.545 3.69 0.545 3.69 0.325 5.82 0.325 5.82 0.61 5.93 0.61 ;
      POLYGON 3.845 0.71 3.485 0.71 3.485 1.09 3.16 1.09 3.16 1.03 3.425 1.03 3.425 0.71 3.16 0.71 3.16 0.455 3.22 0.455 3.22 0.65 3.845 0.65 ;
      POLYGON 3.325 0.93 3.265 0.93 3.265 0.87 3 0.87 3 0.33 2.105 0.33 2.105 0.775 2.135 0.775 2.135 0.835 2.015 0.835 2.015 0.775 2.045 0.775 2.045 0.33 1.755 0.33 1.755 1.02 1.695 1.02 1.695 0.39 1.67 0.39 1.67 0.27 2.28 0.27 2.28 0.215 2.4 0.215 2.4 0.27 3.06 0.27 3.06 0.81 3.325 0.81 ;
      POLYGON 2.9 1.1 2.84 1.1 2.84 0.875 2.45 0.875 2.45 0.815 2.84 0.815 2.84 0.455 2.9 0.455 ;
      POLYGON 2.74 0.715 2.295 0.715 2.295 1.1 2.235 1.1 2.235 0.545 2.205 0.545 2.205 0.485 2.325 0.485 2.325 0.545 2.295 0.545 2.295 0.655 2.74 0.655 ;
      POLYGON 2.04 1.215 0.265 1.215 0.265 1.155 0.64 1.155 0.64 0.59 0.425 0.59 0.425 0.47 0.485 0.47 0.485 0.53 0.7 0.53 0.7 1.155 1.855 1.155 1.855 0.515 1.885 0.515 1.885 0.455 1.945 0.455 1.945 0.575 1.915 0.575 1.915 1.075 2.04 1.075 ;
      POLYGON 1.595 0.695 1.535 0.695 1.535 0.525 1.025 0.525 1.025 0.995 1.385 0.995 1.385 1.055 0.965 1.055 0.965 0.27 1.025 0.27 1.025 0.465 1.595 0.465 ;
  END
END DFFTRX4

MACRO DFFTRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFTRXL 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.29205 LAYER Metal1 ;
    ANTENNADIFFAREA 2.537525 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1944 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.79038075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 90.169753 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.975 0.645 0.94 0.645 0.94 0.9 0.96 0.9 0.96 1.17 0.88 1.17 0.88 0.98 0.86 0.98 0.86 0.57 0.895 0.57 0.895 0.525 0.975 0.525 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.347875 LAYER Metal1 ;
    ANTENNADIFFAREA 2.537525 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1944 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.07754625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 91.37345675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.325 1.02 0.245 1.02 0.245 0.73 0.06 0.73 0.06 0.6 0.245 0.6 0.245 0.54 0.325 0.54 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.37 0.88 4.29 0.88 4.29 0.54 4.26 0.54 4.26 0.41 4.34 0.41 4.34 0.46 4.37 0.46 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.19 0.83 4.06 0.83 4.06 0.38 4.14 0.38 4.14 0.75 4.19 0.75 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 12.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.3 1.01 1.14 1.01 1.14 1.3 1.06 1.3 1.06 0.93 1.22 0.93 1.22 0.89 1.3 0.89 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.77 0 1.77 0 1.65 0.535 1.65 0.535 1.285 0.595 1.285 0.595 1.65 1.07 1.65 1.07 1.51 1.13 1.51 1.13 1.65 1.895 1.65 1.895 1.49 2.015 1.49 2.015 1.55 1.955 1.55 1.955 1.65 2.935 1.65 2.935 1.49 3.055 1.49 3.055 1.55 2.995 1.55 2.995 1.65 4.06 1.65 4.06 1.285 4.12 1.285 4.12 1.65 4.405 1.65 4.405 1.285 4.465 1.285 4.465 1.65 4.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 0.06 4.15 0.06 4.15 0.2 4.09 0.2 4.09 0.06 3.035 0.06 3.035 0.17 2.915 0.17 2.915 0.06 2.01 0.06 2.01 0.63 1.95 0.63 1.95 0.06 1.14 0.06 1.14 0.2 1.08 0.2 1.08 0.06 0.595 0.06 0.595 0.2 0.535 0.2 0.535 0.06 0 0.06 0 -0.06 4.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.53 1.04 4.3 1.04 4.3 1.15 3.57 1.15 3.57 1.21 3.51 1.21 3.51 1.09 3.635 1.09 3.635 0.535 3.695 0.535 3.695 1.09 4.24 1.09 4.24 0.98 4.47 0.98 4.47 0.54 4.53 0.54 ;
      POLYGON 3.915 0.99 3.795 0.99 3.795 0.93 3.855 0.93 3.855 0.435 3.535 0.435 3.535 0.915 3.415 0.915 3.415 0.855 3.475 0.855 3.475 0.435 2.645 0.435 2.645 0.845 2.37 0.845 2.37 0.965 2.31 0.965 2.31 0.785 2.585 0.785 2.585 0.375 3.18 0.375 3.18 0.325 3.3 0.325 3.3 0.375 3.915 0.375 ;
      POLYGON 3.375 0.625 3.315 0.625 3.315 1.015 3.365 1.015 3.365 1.21 3.305 1.21 3.305 1.075 3.255 1.075 3.255 0.945 2.905 0.945 2.905 0.885 3.255 0.885 3.255 0.565 3.375 0.565 ;
      POLYGON 3.33 1.435 3.21 1.435 3.21 1.39 2.58 1.39 2.58 1.435 2.46 1.435 2.46 1.39 1.305 1.39 1.305 1.11 1.4 1.11 1.4 0.54 1.46 0.54 1.46 1.17 1.365 1.17 1.365 1.33 3.27 1.33 3.27 1.375 3.33 1.375 ;
      POLYGON 3.13 0.785 2.805 0.785 2.805 1.18 2.685 1.18 2.685 1.12 2.745 1.12 2.745 0.565 2.865 0.565 2.865 0.725 3.13 0.725 ;
      POLYGON 2.485 0.685 2.21 0.685 2.21 1.12 2.44 1.12 2.44 1.18 2.15 1.18 2.15 1.01 1.79 1.01 1.79 0.95 2.15 0.95 2.15 0.625 2.425 0.625 2.425 0.535 2.485 0.535 ;
      POLYGON 2.05 0.85 1.69 0.85 1.69 1.12 1.78 1.12 1.78 1.18 1.63 1.18 1.63 0.57 1.745 0.57 1.745 0.47 1.56 0.47 1.56 0.44 1.3 0.44 1.3 0.79 1.16 0.79 1.16 0.8 1.04 0.8 1.04 0.73 1.24 0.73 1.24 0.38 1.62 0.38 1.62 0.41 1.805 0.41 1.805 0.63 1.69 0.63 1.69 0.79 1.99 0.79 1.99 0.73 2.05 0.73 ;
      POLYGON 0.76 1.02 0.68 1.02 0.68 0.81 0.425 0.81 0.425 0.73 0.68 0.73 0.68 0.54 0.76 0.54 ;
  END
END DFFTRXL

MACRO DFFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFX1 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.19615 LAYER Metal1 ;
    ANTENNADIFFAREA 2.451875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2205 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.959864 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 76.78911575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 1.34 0.88 1.34 0.88 0.73 0.86 0.73 0.86 0.54 0.94 0.54 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.24795 LAYER Metal1 ;
    ANTENNADIFFAREA 2.451875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2205 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.1947845 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 77.9863945 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.285 1.29 0.205 1.29 0.205 0.73 0.06 0.73 0.06 0.6 0.205 0.6 0.205 0.54 0.285 0.54 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.88 1.085 3.495 1.085 3.495 1.005 3.635 1.005 3.635 0.89 3.715 0.89 3.715 1.005 3.88 1.005 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.285 0.9 1.28 0.9 1.28 1.135 1.06 1.135 1.06 0.98 1.2 0.98 1.2 0.82 1.205 0.82 1.205 0.78 1.285 0.78 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 1.77 0 1.77 0 1.65 0.46 1.65 0.46 1.285 0.52 1.285 0.52 1.65 1.115 1.65 1.115 1.51 1.175 1.51 1.175 1.65 1.79 1.65 1.79 1.54 1.91 1.54 1.91 1.65 2.77 1.65 2.77 1.54 2.89 1.54 2.89 1.65 3.665 1.65 3.665 1.185 3.725 1.185 3.725 1.65 4.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 0.06 3.705 0.06 3.705 0.47 3.645 0.47 3.645 0.06 2.945 0.06 2.945 0.16 3.005 0.16 3.005 0.22 2.885 0.22 2.885 0.06 1.905 0.06 1.905 0.605 1.845 0.605 1.845 0.06 1.125 0.06 1.125 0.52 1.065 0.52 1.065 0.06 0.52 0.06 0.52 0.2 0.46 0.2 0.46 0.06 0 0.06 0 -0.06 4.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.045 0.95 4.04 0.95 4.04 1.21 3.98 1.21 3.98 0.89 3.985 0.89 3.985 0.63 3.465 0.63 3.465 0.41 2.725 0.41 2.725 0.39 2.465 0.39 2.465 0.71 2.53 0.71 2.53 0.83 2.265 0.83 2.265 1.015 2.205 1.015 2.205 0.77 2.405 0.77 2.405 0.33 2.785 0.33 2.785 0.35 3.525 0.35 3.525 0.57 3.88 0.57 3.88 0.51 3.94 0.51 3.94 0.57 4.045 0.57 ;
      POLYGON 3.885 0.79 3.535 0.79 3.535 0.89 3.395 0.89 3.395 1.34 1.385 1.34 1.385 0.54 1.445 0.54 1.445 1.28 2.375 1.28 2.375 0.93 2.435 0.93 2.435 1.28 3.335 1.28 3.335 1.02 3.16 1.02 3.16 0.9 3.22 0.9 3.22 0.96 3.335 0.96 3.335 0.73 3.885 0.73 ;
      POLYGON 3.365 0.63 3.06 0.63 3.06 1.12 3.235 1.12 3.235 1.18 3 1.18 3 0.945 2.85 0.945 2.85 1.005 2.79 1.005 2.79 0.885 3 0.885 3 0.57 3.305 0.57 3.305 0.51 3.365 0.51 ;
      POLYGON 2.9 0.785 2.69 0.785 2.69 1.18 2.535 1.18 2.535 1.12 2.63 1.12 2.63 0.61 2.565 0.61 2.565 0.49 2.625 0.49 2.625 0.55 2.69 0.55 2.69 0.725 2.9 0.725 ;
      POLYGON 2.305 0.6 2.105 0.6 2.105 1.12 2.275 1.12 2.275 1.18 2.045 1.18 2.045 0.985 1.705 0.985 1.705 0.865 1.765 0.865 1.765 0.925 2.045 0.925 2.045 0.54 2.305 0.54 ;
      POLYGON 1.945 0.825 1.885 0.825 1.885 0.765 1.605 0.765 1.605 1.12 1.675 1.12 1.675 1.18 1.545 1.18 1.545 0.545 1.64 0.545 1.64 0.44 1.285 0.44 1.285 0.68 1.1 0.68 1.1 0.82 1.04 0.82 1.04 0.62 1.225 0.62 1.225 0.38 1.7 0.38 1.7 0.605 1.605 0.605 1.605 0.705 1.945 0.705 ;
      POLYGON 0.72 1.02 0.64 1.02 0.64 0.81 0.385 0.81 0.385 0.73 0.64 0.73 0.64 0.54 0.72 0.54 ;
  END
END DFFX1

MACRO DFFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFX2 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5192 LAYER Metal1 ;
    ANTENNADIFFAREA 2.9231 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.285975 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.80916175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 68.051403 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.9 1.29 3.84 1.29 3.84 0.705 3.74 0.705 3.74 0.73 3.66 0.73 3.66 0.6 3.74 0.6 3.74 0.645 3.84 0.645 3.84 0.53 3.9 0.53 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5192 LAYER Metal1 ;
    ANTENNADIFFAREA 2.9231 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.285975 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.80916175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 68.051403 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.53 3.34 1.29 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.86 0.53 2.94 1.03 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.45 1.015 0.365 1.015 0.365 1.275 0.235 1.275 0.235 1.195 0.285 1.195 0.285 0.935 0.37 0.935 0.37 0.895 0.45 0.895 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.305 1.65 0.305 1.375 0.365 1.375 0.365 1.65 1.03 1.65 1.03 1.49 1.15 1.49 1.15 1.55 1.09 1.55 1.09 1.65 2.075 1.65 2.075 1.49 2.195 1.49 2.195 1.55 2.135 1.55 2.135 1.65 3.075 1.65 3.075 1.045 3.135 1.045 3.135 1.65 3.505 1.65 3.505 0.91 3.565 0.91 3.565 1.65 4.045 1.65 4.045 0.93 4.105 0.93 4.105 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 4.22 0.06 4.22 0.51 4.16 0.51 4.16 0.06 3.625 0.06 3.625 0.17 3.505 0.17 3.505 0.06 3.135 0.06 3.135 0.17 3.015 0.17 3.015 0.06 2.195 0.06 2.195 0.575 2.135 0.575 2.135 0.06 1.22 0.06 1.22 0.17 1.1 0.17 1.1 0.06 0.34 0.06 0.34 0.635 0.28 0.635 0.28 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.6 0.62 4.54 0.62 4.54 0.83 4.34 0.83 4.34 1.02 4.28 1.02 4.28 0.83 4 0.83 4 0.77 4.48 0.77 4.48 0.56 4.6 0.56 ;
      POLYGON 4.44 0.425 4.38 0.425 4.38 0.67 4 0.67 4 0.43 3.5 0.43 3.5 0.81 3.44 0.81 3.44 0.43 3.16 0.43 3.16 0.81 3.1 0.81 3.1 0.43 2.4 0.43 2.4 0.53 2.515 0.53 2.515 0.96 2.43 0.96 2.43 1.12 2.31 1.12 2.31 1.06 2.37 1.06 2.37 0.96 2.065 0.96 2.065 0.9 2.455 0.9 2.455 0.59 2.34 0.59 2.34 0.37 4.06 0.37 4.06 0.61 4.32 0.61 4.32 0.365 4.44 0.365 ;
      POLYGON 2.76 1.39 1.665 1.39 1.665 1.4 1.545 1.4 1.545 1.39 0.93 1.39 0.93 1.4 0.755 1.4 0.755 1.34 0.87 1.34 0.87 1.33 2.7 1.33 2.7 0.53 2.76 0.53 ;
      POLYGON 2.355 0.8 2.235 0.8 2.235 0.77 1.965 0.77 1.965 1.15 1.735 1.15 1.735 1.09 1.905 1.09 1.905 0.77 1.64 0.77 1.64 0.54 1.7 0.54 1.7 0.71 2.355 0.71 ;
      POLYGON 1.805 0.99 1.745 0.99 1.745 0.93 1.48 0.93 1.48 0.435 0.61 0.435 0.61 0.86 0.67 0.86 0.67 0.92 0.55 0.92 0.55 0.795 0.13 0.795 0.13 1.175 0.07 1.175 0.07 0.735 0.075 0.735 0.075 0.54 0.135 0.54 0.135 0.735 0.55 0.735 0.55 0.375 0.805 0.375 0.805 0.27 0.925 0.27 0.925 0.375 1.54 0.375 1.54 0.87 1.805 0.87 ;
      POLYGON 1.44 1.145 1.32 1.145 1.32 0.985 0.93 0.985 0.93 0.925 1.32 0.925 1.32 0.535 1.38 0.535 1.38 1.085 1.44 1.085 ;
      POLYGON 1.22 0.8 0.83 0.8 0.83 1.115 0.705 1.115 0.705 1.175 0.645 1.175 0.645 1.055 0.77 1.055 0.77 0.54 0.83 0.54 0.83 0.74 1.22 0.74 ;
  END
END DFFX2

MACRO DFFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFX4 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.081275 LAYER Metal1 ;
    ANTENNADIFFAREA 3.604925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4392 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.0156535 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 54.760929 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.665 0.63 4.14 0.63 4.14 1.015 4.555 1.015 4.555 1.405 4.495 1.405 4.495 1.075 4.145 1.075 4.145 1.405 4.06 1.405 4.06 0.79 4.075 0.79 4.075 0.57 4.665 0.57 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.081275 LAYER Metal1 ;
    ANTENNADIFFAREA 3.604925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4392 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.0156535 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 54.760929 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.735 1.405 3.675 1.405 3.675 1.075 3.325 1.075 3.325 1.405 3.265 1.405 3.265 0.73 3.26 0.73 3.26 0.6 3.28 0.6 3.28 0.5 3.135 0.5 3.135 0.44 3.725 0.44 3.725 0.5 3.34 0.5 3.34 1.015 3.735 1.015 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.525 0.94 1.025 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.24 0.73 0.14 0.73 0.14 0.965 0.06 0.965 0.06 0.565 0.24 0.565 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.065 0.13 1.065 0.13 1.65 0.805 1.65 0.805 1.285 0.865 1.285 0.865 1.65 1.595 1.65 1.595 1.54 1.715 1.54 1.715 1.65 2.62 1.65 2.62 1.095 2.68 1.095 2.68 1.65 3.06 1.65 3.06 1.06 3.12 1.06 3.12 1.65 3.47 1.65 3.47 1.175 3.53 1.175 3.53 1.65 3.88 1.65 3.88 1.015 3.94 1.015 3.94 1.65 4.29 1.65 4.29 1.175 4.35 1.175 4.35 1.65 4.7 1.65 4.7 1.105 4.76 1.105 4.76 1.65 5.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 0.06 4.985 0.06 4.985 0.52 4.925 0.52 4.925 0.06 4.43 0.06 4.43 0.17 4.31 0.17 4.31 0.06 3.96 0.06 3.96 0.17 3.84 0.17 3.84 0.06 3.49 0.06 3.49 0.17 3.37 0.17 3.37 0.06 3.02 0.06 3.02 0.17 2.9 0.17 2.9 0.06 2.52 0.06 2.52 0.2 2.46 0.2 2.46 0.06 1.58 0.06 1.58 0.2 1.52 0.2 1.52 0.06 0.995 0.06 0.995 0.2 0.935 0.2 0.935 0.06 0.13 0.06 0.13 0.465 0.07 0.465 0.07 0.06 0 0.06 0 -0.06 5.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.19 0.68 5.06 0.68 5.06 1.005 4.965 1.005 4.965 1.405 4.905 1.405 4.905 1.005 4.655 1.005 4.655 0.855 4.715 0.855 4.715 0.945 5 0.945 5 0.62 5.13 0.62 5.13 0.54 5.19 0.54 ;
      POLYGON 4.9 0.845 4.84 0.845 4.84 0.755 4.765 0.755 4.765 0.34 2.915 0.34 2.915 0.9 3.1 0.9 3.1 0.84 3.16 0.84 3.16 0.96 2.885 0.96 2.885 1.405 2.825 1.405 2.825 0.96 2.515 0.96 2.515 0.9 2.855 0.9 2.855 0.575 2.695 0.575 2.695 0.455 2.755 0.455 2.755 0.515 2.855 0.515 2.855 0.28 4.825 0.28 4.825 0.695 4.9 0.695 ;
      POLYGON 2.72 0.79 2.255 0.79 2.255 1.22 2.315 1.22 2.315 1.28 2.195 1.28 2.195 0.63 2.16 0.63 2.16 0.57 2.28 0.57 2.28 0.73 2.72 0.73 ;
      POLYGON 2.475 1.44 1.04 1.44 1.04 1.185 0.66 1.185 0.66 1.31 0.57 1.31 0.57 0.605 0.51 0.605 0.51 0.365 0.63 0.365 0.63 1.125 1.04 1.125 1.04 1.02 1.1 1.02 1.1 1.38 2.415 1.38 2.415 1.12 2.355 1.12 2.355 1 2.415 1 2.415 1.06 2.475 1.06 ;
      POLYGON 2.355 0.3 2.295 0.3 2.295 0.36 2.06 0.36 2.06 1.11 2 1.11 2 0.36 1.42 0.36 1.42 1.105 1.36 1.105 1.36 0.36 0.775 0.36 0.775 0.265 0.4 0.265 0.4 1.09 0.34 1.09 0.34 0.205 0.835 0.205 0.835 0.3 1.095 0.3 1.095 0.265 1.215 0.265 1.215 0.3 2.235 0.3 2.235 0.24 2.355 0.24 ;
      POLYGON 2.095 1.28 1.975 1.28 1.975 1.27 1.84 1.27 1.84 0.845 1.53 0.845 1.53 0.725 1.59 0.725 1.59 0.785 1.84 0.785 1.84 0.54 1.9 0.54 1.9 1.21 2.035 1.21 2.035 1.22 2.095 1.22 ;
      POLYGON 1.74 1.095 1.58 1.095 1.58 1.265 1.32 1.265 1.32 1.28 1.2 1.28 1.2 0.63 1.14 0.63 1.14 0.57 1.26 0.57 1.26 1.205 1.52 1.205 1.52 1.035 1.74 1.035 ;
  END
END DFFX4

MACRO DFFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFXL 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5502 LAYER Metal1 ;
    ANTENNADIFFAREA 2.27205 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1944 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.11831275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 102.06790125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.055 1.115 0.94 1.115 0.94 1.3 0.86 1.3 0.86 0.56 0.92 0.56 0.92 0.52 1 0.52 1 0.64 0.94 0.64 0.94 0.995 1.055 0.995 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5502 LAYER Metal1 ;
    ANTENNADIFFAREA 2.27205 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1944 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.11831275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 102.06790125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.35 0.66 0.27 0.66 0.27 0.94 0.35 0.94 0.35 1.06 0.27 1.06 0.27 1.02 0.19 1.02 0.19 0.73 0.06 0.73 0.06 0.54 0.35 0.54 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.17 1.085 4.14 1.085 4.14 1.185 3.93 1.185 3.93 0.845 4.17 0.845 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.565 0.895 1.3 0.895 1.3 0.79 1.26 0.79 1.26 0.62 1.38 0.62 1.38 0.815 1.565 0.815 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.495 1.65 0.495 0.995 0.555 0.995 0.555 1.65 1.2 1.65 1.2 0.995 1.26 0.995 1.26 1.65 2.06 1.65 2.06 1.54 2.18 1.54 2.18 1.65 3.13 1.65 3.13 1.54 3.25 1.54 3.25 1.65 4.045 1.65 4.045 1.285 4.105 1.285 4.105 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 4.105 0.06 4.105 0.365 3.985 0.365 3.985 0.305 4.045 0.305 4.045 0.06 3.35 0.06 3.35 0.25 3.23 0.25 3.23 0.19 3.29 0.19 3.29 0.06 2.105 0.06 2.105 0.43 2.045 0.43 2.045 0.06 1.165 0.06 1.165 0.2 1.105 0.2 1.105 0.06 0.555 0.06 0.555 0.635 0.495 0.635 0.495 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.33 1.31 4.27 1.31 4.27 0.525 3.825 0.525 3.825 0.235 3.51 0.235 3.51 0.41 3.07 0.41 3.07 0.235 2.81 0.235 2.81 0.685 2.45 0.685 2.45 1.02 2.39 1.02 2.39 0.625 2.75 0.625 2.75 0.175 3.13 0.175 3.13 0.35 3.45 0.35 3.45 0.175 3.885 0.175 3.885 0.465 4.25 0.465 4.25 0.335 4.33 0.335 ;
      POLYGON 4.17 0.745 3.83 0.745 3.83 1.47 3.33 1.47 3.33 1.44 2.75 1.44 2.75 1.47 2.37 1.47 2.37 1.44 1.43 1.44 1.43 0.995 1.665 0.995 1.665 0.635 1.545 0.635 1.545 0.515 1.605 0.515 1.605 0.575 1.725 0.575 1.725 1.055 1.49 1.055 1.49 1.38 2.43 1.38 2.43 1.41 2.69 1.41 2.69 1.06 2.81 1.06 2.81 1.12 2.75 1.12 2.75 1.38 3.39 1.38 3.39 1.41 3.77 1.41 3.77 1.035 3.49 1.035 3.49 0.975 3.77 0.975 3.77 0.685 3.805 0.685 3.805 0.625 3.865 0.625 3.865 0.685 4.17 0.685 ;
      POLYGON 3.725 0.455 3.67 0.455 3.67 0.8 3.39 0.8 3.39 1.135 3.62 1.135 3.62 1.31 3.56 1.31 3.56 1.195 3.33 1.195 3.33 0.8 3.13 0.8 3.13 0.86 3.07 0.86 3.07 0.74 3.61 0.74 3.61 0.395 3.665 0.395 3.665 0.335 3.725 0.335 ;
      POLYGON 3.23 0.64 2.97 0.64 2.97 1.28 2.85 1.28 2.85 1.22 2.91 1.22 2.91 0.335 2.97 0.335 2.97 0.58 3.17 0.58 3.17 0.52 3.23 0.52 ;
      POLYGON 2.65 0.425 2.29 0.425 2.29 1.12 2.59 1.12 2.59 1.31 2.53 1.31 2.53 1.18 2.23 1.18 2.23 0.87 2.045 0.87 2.045 0.75 2.105 0.75 2.105 0.81 2.23 0.81 2.23 0.365 2.65 0.365 ;
      POLYGON 2.13 0.65 1.945 0.65 1.945 1.28 1.825 1.28 1.825 1.22 1.885 1.22 1.885 0.65 1.825 0.65 1.825 0.395 1.325 0.395 1.325 0.52 1.16 0.52 1.16 0.8 1.04 0.8 1.04 0.74 1.1 0.74 1.1 0.46 1.265 0.46 1.265 0.335 1.885 0.335 1.885 0.59 2.07 0.59 2.07 0.53 2.13 0.53 ;
      POLYGON 0.76 1.02 0.68 1.02 0.68 0.84 0.4 0.84 0.4 0.76 0.68 0.76 0.68 0.54 0.76 0.54 ;
  END
END DFFXL

MACRO DLY1X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY1X1 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9033 LAYER Metal1 ;
    ANTENNADIFFAREA 0.9218 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.07785 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.60308275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 94.79768775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.52 1.74 1.29 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 0.94 0.46 0.94 0.46 0.895 0.28 0.895 0.28 0.775 0.46 0.775 0.46 0.62 0.54 0.62 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.355 1.65 0.355 1.04 0.415 1.04 0.415 1.65 0.64 1.65 0.64 0.63 0.76 0.63 0.76 0.69 0.7 0.69 0.7 1.65 1.455 1.65 1.455 1.08 1.515 1.08 1.515 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.515 0.06 1.515 0.5 1.455 0.5 1.455 0.06 0.7 0.06 0.7 0.47 0.92 0.47 0.92 0.85 0.8 0.85 0.8 0.79 0.86 0.79 0.86 0.53 0.64 0.53 0.64 0.06 0.415 0.06 0.415 0.355 0.355 0.355 0.355 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.56 0.98 1.28 0.98 1.28 1.04 1.22 1.04 1.22 0.92 1.5 0.92 1.5 0.66 1.22 0.66 1.22 0.52 1.28 0.52 1.28 0.6 1.56 0.6 ;
      POLYGON 1.385 0.82 1.08 0.82 1.08 1.01 0.86 1.01 0.86 1.07 0.8 1.07 0.8 0.95 1.02 0.95 1.02 0.37 0.8 0.37 0.8 0.25 0.86 0.25 0.86 0.31 1.08 0.31 1.08 0.76 1.385 0.76 ;
      POLYGON 0.52 0.52 0.18 0.52 0.18 1.065 0.12 1.065 0.12 0.26 0.18 0.26 0.18 0.46 0.52 0.46 ;
  END
END DLY1X1

MACRO DLY1X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY1X4 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2673 LAYER Metal1 ;
    ANTENNADIFFAREA 1.322975 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.17865 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.09375875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 57.6490345 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.905 0.66 1.52 0.66 1.52 0.79 1.54 0.79 1.54 0.9 1.905 0.9 1.905 1.29 1.845 1.29 1.845 0.96 1.495 0.96 1.495 1.29 1.435 1.29 1.435 0.9 1.46 0.9 1.46 0.66 1.435 0.66 1.435 0.52 1.495 0.52 1.495 0.6 1.845 0.6 1.845 0.52 1.905 0.52 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.445 0.895 0.315 0.895 0.315 1.145 0.235 1.145 0.235 0.775 0.445 0.775 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.37 1.65 0.37 1.245 0.43 1.245 0.43 1.65 0.545 1.65 0.545 0.775 0.605 0.775 0.605 1.65 1.23 1.65 1.23 1.08 1.29 1.08 1.29 1.65 1.64 1.65 1.64 1.06 1.7 1.06 1.7 1.65 2.05 1.65 2.05 0.9 2.11 0.9 2.11 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 2.11 0.06 2.11 0.5 2.05 0.5 2.05 0.06 1.7 0.06 1.7 0.5 1.64 0.5 1.64 0.06 1.29 0.06 1.29 0.5 1.23 0.5 1.23 0.06 0.605 0.06 0.605 0.615 0.765 0.615 0.765 1.075 0.705 1.075 0.705 0.675 0.545 0.675 0.545 0.06 0.375 0.06 0.375 0.515 0.315 0.515 0.315 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.335 0.98 1.085 0.98 1.085 1.29 1.025 1.29 1.025 0.92 1.275 0.92 1.275 0.66 1.025 0.66 1.025 0.52 1.085 0.52 1.085 0.6 1.335 0.6 ;
      POLYGON 1.175 0.82 0.925 0.82 0.925 1.235 0.765 1.235 0.765 1.295 0.705 1.295 0.705 1.175 0.865 1.175 0.865 0.515 0.705 0.515 0.705 0.395 0.765 0.395 0.765 0.455 0.925 0.455 0.925 0.76 1.175 0.76 ;
      POLYGON 0.445 0.675 0.135 0.675 0.135 1.245 0.225 1.245 0.225 1.365 0.165 1.365 0.165 1.305 0.075 1.305 0.075 0.455 0.11 0.455 0.11 0.395 0.17 0.395 0.17 0.515 0.135 0.515 0.135 0.615 0.445 0.615 ;
  END
END DLY1X4

MACRO DLY2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY2X1 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.997775 LAYER Metal1 ;
    ANTENNADIFFAREA 1.70205 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.14265 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.00473175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 114.7423765 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.33 0.475 0.14 0.475 0.14 1.115 0.33 1.115 0.33 1.395 0.27 1.395 0.27 1.175 0.08 1.175 0.08 0.73 0.06 0.73 0.06 0.6 0.08 0.6 0.08 0.415 0.27 0.415 0.27 0.355 0.33 0.355 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 0.73 1.52 0.73 1.52 1.08 1.44 1.08 1.44 0.625 1.46 0.625 1.46 0.6 1.54 0.6 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 1.77 0 1.77 0 1.65 0.43 1.65 0.43 1.015 0.24 1.015 0.24 0.575 0.82 0.575 0.82 0.635 0.3 0.635 0.3 0.955 0.49 0.955 0.49 1.275 0.535 1.275 0.535 1.65 1.485 1.65 1.485 1.49 1.605 1.49 1.605 1.55 1.545 1.55 1.545 1.65 2.65 1.65 2.65 1.23 2.355 1.23 2.355 0.725 2.415 0.725 2.415 0.85 2.985 0.85 2.985 0.91 2.415 0.91 2.415 1.17 2.71 1.17 2.71 1.65 3.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 0.06 3.115 0.06 3.115 0.69 3.145 0.69 3.145 1.13 2.97 1.13 2.97 1.01 3.085 1.01 3.085 0.75 3.055 0.75 3.055 0.06 2.735 0.06 2.735 0.5 2.795 0.5 2.795 0.56 2.675 0.56 2.675 0.06 1.935 0.06 1.935 0.6 1.85 0.6 1.85 0.95 1.79 0.95 1.79 0.54 1.875 0.54 1.875 0.06 1.535 0.06 1.535 0.17 1.415 0.17 1.415 0.06 0.98 0.06 0.98 0.855 0.92 0.855 0.92 0.06 0.535 0.06 0.535 0.475 0.475 0.475 0.475 0.06 0 0.06 0 -0.06 3.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.305 1.295 2.81 1.295 2.81 1.07 2.555 1.07 2.555 1.01 2.87 1.01 2.87 1.235 3.245 1.235 3.245 0.59 3.215 0.59 3.215 0.47 3.275 0.47 3.275 0.53 3.305 0.53 ;
      POLYGON 2.955 0.72 2.515 0.72 2.515 0.395 2.095 0.395 2.095 1.11 1.915 1.11 1.915 1.17 1.855 1.17 1.855 1.05 2.035 1.05 2.035 0.335 2.575 0.335 2.575 0.66 2.895 0.66 2.895 0.4 2.835 0.4 2.835 0.34 2.955 0.34 ;
      POLYGON 2.535 1.39 1.385 1.39 1.385 1.445 0.635 1.445 0.635 1.175 0.59 1.175 0.59 0.855 0.4 0.855 0.4 0.735 0.46 0.735 0.46 0.795 0.65 0.795 0.65 1.115 0.695 1.115 0.695 1.385 1.325 1.385 1.325 1.33 2.195 1.33 2.195 0.565 2.355 0.565 2.355 0.495 2.415 0.495 2.415 0.625 2.255 0.625 2.255 1.33 2.535 1.33 ;
      POLYGON 1.775 0.44 1.14 0.44 1.14 1.065 1.045 1.065 1.045 1.125 0.985 1.125 0.985 1.005 1.08 1.005 1.08 0.38 1.775 0.38 ;
      POLYGON 1.34 1.23 1.225 1.23 1.225 1.285 0.795 1.285 0.795 1.015 0.75 1.015 0.75 0.835 0.81 0.835 0.81 0.955 0.855 0.955 0.855 1.225 1.165 1.225 1.165 1.17 1.28 1.17 1.28 0.54 1.34 0.54 ;
  END
END DLY2X1

MACRO DLY2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY2X4 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.14 1.075 2.035 1.075 2.035 0.84 2.06 0.84 2.06 0.6 2.14 0.6 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.34175 LAYER Metal1 ;
    ANTENNADIFFAREA 2.321525 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.24345 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.61901825 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 76.66050525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.835 0.475 0.79 0.475 0.79 1.115 0.835 1.115 0.835 1.335 0.775 1.335 0.775 1.175 0.73 1.175 0.73 0.66 0.54 0.66 0.54 0.73 0.425 0.73 0.425 1.335 0.365 1.335 0.365 0.495 0.425 0.495 0.425 0.6 0.73 0.6 0.73 0.415 0.775 0.415 0.775 0.355 0.835 0.355 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 0 1.77 0 1.65 0.16 1.65 0.16 0.945 0.22 0.945 0.22 1.65 0.57 1.65 0.57 0.945 0.63 0.945 0.63 1.65 0.935 1.65 0.935 1.015 0.89 1.015 0.89 0.575 1.415 0.575 1.415 0.635 0.95 0.635 0.95 0.955 0.995 0.955 0.995 1.215 1.04 1.215 1.04 1.335 0.995 1.335 0.995 1.65 2.11 1.65 2.11 1.51 2.17 1.51 2.17 1.65 3.01 1.65 3.01 0.815 2.95 0.815 2.95 0.755 3.07 0.755 3.07 0.78 3.61 0.78 3.61 0.84 3.07 0.84 3.07 1.65 4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.77 0.06 3.77 1.06 3.52 1.06 3.52 0.94 3.71 0.94 3.71 0.06 3.39 0.06 3.39 0.43 3.45 0.43 3.45 0.49 3.33 0.49 3.33 0.06 2.53 0.06 2.53 0.93 2.345 0.93 2.345 0.87 2.47 0.87 2.47 0.06 2.13 0.06 2.13 0.17 2.01 0.17 2.01 0.06 1.575 0.06 1.575 0.795 1.415 0.795 1.415 0.735 1.515 0.735 1.515 0.06 1.14 0.06 1.14 0.475 1.08 0.475 1.08 0.06 0.63 0.06 0.63 0.475 0.57 0.475 0.57 0.06 0.22 0.06 0.22 0.475 0.16 0.475 0.16 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.93 1.22 3.17 1.22 3.17 0.94 3.23 0.94 3.23 1.16 3.87 1.16 3.87 0.4 3.93 0.4 ;
      POLYGON 3.61 0.65 3.17 0.65 3.17 0.47 2.69 0.47 2.69 1.09 2.51 1.09 2.51 1.15 2.45 1.15 2.45 1.03 2.63 1.03 2.63 0.41 3.23 0.41 3.23 0.59 3.55 0.59 3.55 0.33 3.49 0.33 3.49 0.27 3.61 0.27 ;
      POLYGON 3.07 0.63 2.85 0.63 2.85 1.07 2.865 1.07 2.865 1.46 2.805 1.46 2.805 1.31 2.01 1.31 2.01 1.355 1.14 1.355 1.14 1.115 1.095 1.115 1.095 0.855 1.05 0.855 1.05 0.735 1.11 0.735 1.11 0.795 1.155 0.795 1.155 1.055 1.2 1.055 1.2 1.295 1.95 1.295 1.95 1.25 2.79 1.25 2.79 0.57 3.07 0.57 ;
      POLYGON 2.37 0.44 1.735 0.44 1.735 0.99 1.58 0.99 1.58 1.035 1.46 1.035 1.46 0.975 1.52 0.975 1.52 0.93 1.675 0.93 1.675 0.38 2.37 0.38 ;
      POLYGON 1.935 1.15 1.74 1.15 1.74 1.195 1.3 1.195 1.3 0.955 1.255 0.955 1.255 0.775 1.315 0.775 1.315 0.895 1.36 0.895 1.36 1.135 1.68 1.135 1.68 1.09 1.875 1.09 1.875 0.54 1.935 0.54 ;
  END
END DLY2X4

MACRO DLY3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY3X1 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7696 LAYER Metal1 ;
    ANTENNADIFFAREA 2.36775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20745 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.350687 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 108.6550975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.89 1.29 2.83 1.29 2.83 0.895 2.635 0.895 2.635 0.54 2.695 0.54 2.695 0.815 2.89 0.815 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.935 1.065 1.66 1.065 1.66 0.79 1.755 0.79 1.755 0.76 1.935 0.76 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.785 1.65 0.785 1.165 0.7 1.165 0.7 1.105 0.845 1.105 0.845 1.18 0.96 1.18 0.96 0.685 0.455 0.685 0.455 0.625 1.08 0.625 1.08 0.685 1.02 0.685 1.02 1.24 0.845 1.24 0.845 1.65 1.82 1.65 1.82 1.165 1.88 1.165 1.88 1.65 2.035 1.65 2.035 0.76 2.155 0.76 2.155 0.82 2.095 0.82 2.095 1.65 3.065 1.65 3.065 1.26 3.005 1.26 3.005 1.2 3.125 1.2 3.125 1.65 3.875 1.65 3.875 0.7 4.45 0.7 4.45 0.76 3.935 0.76 3.935 1.65 4.115 1.65 4.115 1.115 4.175 1.115 4.175 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 4.53 0.06 4.53 0.54 4.61 0.54 4.61 0.98 4.435 0.98 4.435 0.86 4.55 0.86 4.55 0.6 4.47 0.6 4.47 0.06 4.15 0.06 4.15 0.32 4.21 0.32 4.21 0.44 4.15 0.44 4.15 0.38 4.09 0.38 4.09 0.06 3.455 0.06 3.455 0.81 3.29 0.81 3.29 0.75 3.395 0.75 3.395 0.06 3.075 0.06 3.075 0.49 2.955 0.49 2.955 0.43 3.015 0.43 3.015 0.06 2.315 0.06 2.315 0.915 2.375 0.915 2.375 0.975 2.255 0.975 2.255 0.06 1.88 0.06 1.88 0.5 1.82 0.5 1.82 0.06 1.2 0.06 1.2 0.465 1.24 0.465 1.24 0.82 1.18 0.82 1.18 0.525 1.14 0.525 1.14 0.06 0.79 0.06 0.79 0.365 0.73 0.365 0.73 0.06 0.355 0.06 0.355 0.785 0.575 0.785 0.575 0.845 0.295 0.845 0.295 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.77 1.14 4.275 1.14 4.275 0.925 4.035 0.925 4.035 0.865 4.335 0.865 4.335 1.08 4.71 1.08 4.71 0.44 4.63 0.44 4.63 0.32 4.69 0.32 4.69 0.38 4.77 0.38 ;
      POLYGON 4.37 0.6 3.93 0.6 3.93 0.245 3.615 0.245 3.615 0.97 3.445 0.97 3.445 1.03 3.385 1.03 3.385 0.91 3.555 0.91 3.555 0.185 3.99 0.185 3.99 0.54 4.31 0.54 4.31 0.22 4.25 0.22 4.25 0.16 4.37 0.16 ;
      POLYGON 3.83 0.465 3.775 0.465 3.775 1.19 3.225 1.19 3.225 1.1 3.13 1.1 3.13 0.83 2.99 0.83 2.99 0.77 3.19 0.77 3.19 1.04 3.285 1.04 3.285 1.13 3.715 1.13 3.715 0.405 3.77 0.405 3.77 0.345 3.83 0.345 ;
      POLYGON 3.295 0.335 3.235 0.335 3.235 0.65 2.795 0.65 2.795 0.44 2.475 0.44 2.475 0.54 2.535 0.54 2.535 1.135 2.255 1.135 2.255 1.195 2.195 1.195 2.195 1.075 2.475 1.075 2.475 0.6 2.415 0.6 2.415 0.38 2.855 0.38 2.855 0.59 3.175 0.59 3.175 0.275 3.295 0.275 ;
      POLYGON 2.1 0.31 2.04 0.31 2.04 0.66 1.66 0.66 1.66 0.305 1.4 0.305 1.4 1.1 1.34 1.1 1.34 0.365 1.3 0.365 1.3 0.245 1.72 0.245 1.72 0.6 1.98 0.6 1.98 0.25 2.1 0.25 ;
      POLYGON 1.675 1.4 0.945 1.4 0.945 1.34 1.615 1.34 1.615 1.225 1.5 1.225 1.5 0.405 1.56 0.405 1.56 1.165 1.675 1.165 ;
      POLYGON 0.86 0.91 0.735 0.91 0.735 1.005 0.48 1.005 0.48 1.1 0.42 1.1 0.42 1.005 0.135 1.005 0.135 0.27 0.195 0.27 0.195 0.945 0.675 0.945 0.675 0.85 0.86 0.85 ;
  END
END DLY3X1

MACRO DLY3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY3X4 0 0 ;
  SIZE 5.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 0.73 1.66 0.73 1.66 1.02 1.58 1.02 1.58 0.61 1.66 0.61 1.66 0.6 1.74 0.6 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.05195 LAYER Metal1 ;
    ANTENNADIFFAREA 2.93975 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.30825 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.90089225 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 77.76155725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.03 0.535 3.01 0.535 3.01 1.29 2.95 1.29 2.95 0.66 2.6 0.66 2.6 1.29 2.54 1.29 2.54 0.73 2.46 0.73 2.46 0.535 2.44 0.535 2.44 0.475 2.56 0.475 2.56 0.6 2.91 0.6 2.91 0.475 3.03 0.475 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.2 1.77 0 1.77 0 1.65 0.645 1.65 0.645 1.18 0.56 1.18 0.56 1.12 0.645 1.12 0.645 1.025 0.82 1.025 0.82 0.765 0.415 0.765 0.415 0.6 0.535 0.6 0.535 0.705 0.94 0.705 0.94 0.765 0.88 0.765 0.88 1.085 0.705 1.085 0.705 1.65 1.625 1.65 1.625 1.12 1.685 1.12 1.685 1.65 1.84 1.65 1.84 0.895 1.96 0.895 1.96 0.955 1.9 0.955 1.9 1.65 2.335 1.65 2.335 1.17 2.395 1.17 2.395 1.65 2.745 1.65 2.745 0.9 2.805 0.9 2.805 1.65 3.155 1.65 3.155 1.06 3.215 1.06 3.215 1.65 4.26 1.65 4.26 0.72 4.15 0.72 4.15 0.66 4.795 0.66 4.795 0.78 4.735 0.78 4.735 0.72 4.32 0.72 4.32 1.65 5.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.2 0.06 4.895 0.06 4.895 0.5 4.955 0.5 4.955 0.95 4.895 0.95 4.895 0.56 4.835 0.56 4.835 0.06 4.515 0.06 4.515 0.4 4.395 0.4 4.395 0.34 4.455 0.34 4.455 0.06 3.73 0.06 3.73 0.89 3.66 0.89 3.66 0.77 3.67 0.77 3.67 0.06 3.35 0.06 3.35 0.45 3.41 0.45 3.41 0.51 3.29 0.51 3.29 0.06 2.795 0.06 2.795 0.17 2.675 0.17 2.675 0.06 2.18 0.06 2.18 0.2 2.12 0.2 2.12 0.06 2.005 0.06 2.005 0.735 2.12 0.735 2.12 0.865 2.06 0.865 2.06 0.795 1.945 0.795 1.945 0.06 1.675 0.06 1.675 0.17 1.555 0.17 1.555 0.06 0.91 0.06 0.91 0.545 1.1 0.545 1.1 0.925 0.98 0.925 0.98 0.865 1.04 0.865 1.04 0.605 0.85 0.605 0.85 0.06 0.75 0.06 0.75 0.445 0.69 0.445 0.69 0.06 0.315 0.06 0.315 0.86 0.255 0.86 0.255 0.06 0 0.06 0 -0.06 5.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.115 1.115 4.735 1.115 4.735 0.94 4.42 0.94 4.42 0.82 4.54 0.82 4.54 0.88 4.795 0.88 4.795 1.055 5.055 1.055 5.055 0.4 4.995 0.4 4.995 0.34 5.115 0.34 ;
      POLYGON 4.735 0.24 4.675 0.24 4.675 0.56 4.235 0.56 4.235 0.38 3.89 0.38 3.89 1.05 3.71 1.05 3.71 1.11 3.65 1.11 3.65 0.99 3.83 0.99 3.83 0.32 4.295 0.32 4.295 0.5 4.615 0.5 4.615 0.18 4.735 0.18 ;
      POLYGON 4.135 0.54 4.05 0.54 4.05 0.92 4.115 0.92 4.115 1.31 4.055 1.31 4.055 1.27 3.315 1.27 3.315 0.83 3.11 0.83 3.11 0.77 3.375 0.77 3.375 1.21 3.99 1.21 3.99 0.48 4.135 0.48 ;
      POLYGON 3.57 0.67 3.13 0.67 3.13 0.375 2.34 0.375 2.34 0.575 2.28 0.575 2.28 1.025 2.195 1.025 2.195 1.145 2.135 1.145 2.135 0.965 2.22 0.965 2.22 0.635 2.105 0.635 2.105 0.515 2.28 0.515 2.28 0.315 3.19 0.315 3.19 0.61 3.51 0.61 3.51 0.35 3.45 0.35 3.45 0.29 3.57 0.29 ;
      POLYGON 1.845 0.445 1.26 0.445 1.26 1.085 1.21 1.085 1.21 1.145 1.15 1.145 1.15 1.025 1.2 1.025 1.2 0.445 1.01 0.445 1.01 0.325 1.07 0.325 1.07 0.385 1.845 0.385 ;
      POLYGON 1.48 1.415 0.805 1.415 0.805 1.355 1.42 1.355 1.42 0.63 1.36 0.63 1.36 0.57 1.48 0.57 ;
      POLYGON 0.72 0.925 0.545 0.925 0.545 1.02 0.295 1.02 0.295 1.085 0.095 1.085 0.095 0.35 0.155 0.35 0.155 0.96 0.485 0.96 0.485 0.865 0.72 0.865 ;
  END
END DLY3X4

MACRO DLY4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY4X1 0 0 ;
  SIZE 5.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.2709 LAYER Metal1 ;
    ANTENNADIFFAREA 3.016875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.27225 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.014325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 94.04958675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.565 0.705 0.515 0.705 0.515 1.29 0.435 1.29 0.435 0.54 0.515 0.54 0.515 0.625 0.565 0.625 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.46 0.69 5.54 1.19 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 1.77 0 1.77 0 1.65 0.23 1.65 0.23 0.9 0.29 0.9 0.29 1.65 0.825 1.65 0.825 0.715 1.39 0.715 1.39 0.775 0.885 0.775 0.885 1.54 1.095 1.54 1.095 1.65 1.81 1.65 1.81 1.415 1.75 1.415 1.75 1.355 1.87 1.355 1.87 1.65 2.405 1.65 2.405 0.765 2.345 0.765 2.345 0.705 2.465 0.705 2.465 1.65 3.055 1.65 3.055 1.54 3.175 1.54 3.175 1.65 4.215 1.65 4.215 0.74 4.155 0.74 4.155 0.665 4.74 0.665 4.74 0.785 4.68 0.785 4.68 0.725 4.275 0.725 4.275 1.65 4.485 1.65 4.485 1.51 4.545 1.51 4.545 1.65 5.435 1.65 5.435 1.29 5.495 1.29 5.495 1.65 5.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 0.06 5.495 0.06 5.495 0.425 5.435 0.425 5.435 0.06 5.26 0.06 5.26 0.71 5.25 0.71 5.25 0.94 5.19 0.94 5.19 0.65 5.2 0.65 5.2 0.06 4.455 0.06 4.455 0.2 4.395 0.2 4.395 0.06 4.055 0.06 4.055 0.91 3.935 0.91 3.935 0.85 3.995 0.85 3.995 0.06 3.515 0.06 3.515 0.87 3.395 0.87 3.395 0.81 3.455 0.81 3.455 0.06 3.02 0.06 3.02 0.2 2.96 0.2 2.96 0.06 2.625 0.06 2.625 1.1 2.565 1.1 2.565 0.06 2.075 0.06 2.075 1.025 2.145 1.025 2.145 1.085 2.015 1.085 2.015 0.06 1.84 0.06 1.84 0.2 1.78 0.2 1.78 0.06 1.55 0.06 1.55 0.93 1.49 0.93 1.49 0.06 1.115 0.06 1.115 0.615 1.055 0.615 1.055 0.06 0.175 0.06 0.175 0.52 0.115 0.52 0.115 0.06 0 0.06 0 -0.06 5.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.7 1.36 5.64 1.36 5.64 0.59 5.36 0.59 5.36 0.53 5.64 0.53 5.64 0.33 5.7 0.33 ;
      POLYGON 5.185 1.315 5.125 1.315 5.125 1.255 5.03 1.255 5.03 0.49 5.04 0.49 5.04 0.39 4.555 0.39 4.555 0.33 5.1 0.33 5.1 0.55 5.09 0.55 5.09 1.195 5.185 1.195 ;
      POLYGON 4.9 0.945 4.815 0.945 4.815 1.125 4.755 1.125 4.755 0.945 4.375 0.945 4.375 0.875 4.495 0.875 4.495 0.885 4.84 0.885 4.84 0.49 4.9 0.49 ;
      POLYGON 4.115 1.19 3.065 1.19 3.065 0.3 3.12 0.3 3.12 0.16 3.24 0.16 3.24 0.36 3.125 0.36 3.125 1.13 3.775 1.13 3.775 0.55 3.835 0.55 3.835 0.49 3.895 0.49 3.895 0.61 3.835 0.61 3.835 1.13 4.115 1.13 ;
      POLYGON 3.675 1.03 3.225 1.03 3.225 0.97 3.615 0.97 3.615 0.49 3.675 0.49 ;
      POLYGON 3.58 1.35 2.905 1.35 2.905 0.72 2.8 0.72 2.8 0.32 2.725 0.32 2.725 0.26 2.86 0.26 2.86 0.66 2.965 0.66 2.965 1.29 3.58 1.29 ;
      RECT 2.725 0.82 2.805 1.32 ;
      POLYGON 2.465 0.56 2.345 0.56 2.345 0.34 2.185 0.34 2.185 0.26 2.425 0.26 2.425 0.48 2.465 0.48 ;
      POLYGON 2.305 1.255 2.18 1.255 2.18 1.315 2.12 1.315 2.12 1.255 1.265 1.255 1.265 1.35 1.145 1.35 1.145 1.29 1.205 1.29 1.205 1.195 2.245 1.195 2.245 0.925 2.175 0.925 2.175 0.49 2.235 0.49 2.235 0.865 2.305 0.865 ;
      POLYGON 1.71 1.095 1.33 1.095 1.33 0.935 0.985 0.935 0.985 0.875 1.39 0.875 1.39 1.035 1.65 1.035 1.65 0.52 1.71 0.52 ;
      POLYGON 0.91 0.615 0.725 0.615 0.725 1.125 0.665 1.125 0.665 0.555 0.85 0.555 0.85 0.44 0.335 0.44 0.335 0.79 0.215 0.79 0.215 0.73 0.275 0.73 0.275 0.38 0.91 0.38 ;
  END
END DLY4X1

MACRO DLY4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DLY4X4 0 0 ;
  SIZE 6.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.97 1.06 5.94 1.06 5.94 1.235 5.86 1.235 5.86 0.98 5.89 0.98 5.89 0.765 5.97 0.765 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.423 LAYER Metal1 ;
    ANTENNADIFFAREA 3.4161 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.37305 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.17571375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 71.5641335 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.16 0.99 1.04 0.99 1.04 0.93 1.07 0.93 1.07 0.73 0.72 0.73 0.72 0.99 0.57 0.99 0.57 0.93 0.66 0.93 0.66 0.49 0.72 0.49 0.72 0.6 0.74 0.6 0.74 0.67 1.07 0.67 1.07 0.49 1.13 0.49 1.13 0.93 1.16 0.93 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 0 1.77 0 1.65 0.31 1.65 0.31 1.25 0.43 1.25 0.43 1.31 0.37 1.31 0.37 1.65 0.805 1.65 0.805 1.25 0.925 1.25 0.925 1.31 0.865 1.31 0.865 1.65 1.305 1.65 1.305 1.25 1.365 1.25 1.365 1.65 1.875 1.65 1.875 1.395 1.995 1.395 1.995 1.455 1.935 1.455 1.935 1.65 2.69 1.65 2.69 1.05 2.75 1.05 2.75 1.65 3.48 1.65 3.48 1.55 3.42 1.55 3.42 1.49 3.54 1.49 3.54 1.65 4.51 1.65 4.51 0.715 4.5 0.715 4.5 0.595 5.1 0.595 5.1 0.72 5.04 0.72 5.04 0.655 4.57 0.655 4.57 1.65 4.735 1.65 4.735 1.01 4.795 1.01 4.795 1.65 5.835 1.65 5.835 1.51 5.895 1.51 5.895 1.65 6.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 5.885 0.06 5.885 0.5 5.825 0.5 5.825 0.06 5.62 0.06 5.62 0.85 5.56 0.85 5.56 0.06 4.825 0.06 4.825 0.2 4.765 0.2 4.765 0.06 4.4 0.06 4.4 0.77 4.39 0.77 4.39 0.83 4.33 0.83 4.33 0.71 4.34 0.71 4.34 0.06 3.88 0.06 3.88 0.78 3.76 0.78 3.76 0.72 3.82 0.72 3.82 0.06 3.49 0.06 3.49 0.46 3.43 0.46 3.43 0.06 2.93 0.06 2.93 0.89 2.99 0.89 2.99 0.95 2.87 0.95 2.87 0.06 2.37 0.06 2.37 0.565 2.43 0.565 2.43 1.045 2.18 1.045 2.18 0.925 2.37 0.925 2.37 0.625 2.31 0.625 2.31 0.06 2.21 0.06 2.21 0.495 2.15 0.495 2.15 0.06 1.575 0.06 1.575 0.675 1.635 0.675 1.635 0.795 1.575 0.795 1.575 0.735 1.515 0.735 1.515 0.06 1.335 0.06 1.335 0.47 1.275 0.47 1.275 0.06 0.925 0.06 0.925 0.47 0.865 0.47 0.865 0.06 0.515 0.06 0.515 0.47 0.455 0.47 0.455 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.13 1.055 6.07 1.055 6.07 0.665 5.72 0.665 5.72 0.605 6.03 0.605 6.03 0.405 6.09 0.405 6.09 0.605 6.13 0.605 ;
      POLYGON 5.555 1.07 5.495 1.07 5.495 1.01 5.4 1.01 5.4 0.325 4.925 0.325 4.925 0.265 5.46 0.265 5.46 0.95 5.555 0.95 ;
      POLYGON 5.26 0.88 5.175 0.88 5.175 1.035 5.115 1.035 5.115 0.88 4.67 0.88 4.67 0.755 4.73 0.755 4.73 0.82 5.2 0.82 5.2 0.425 5.26 0.425 ;
      POLYGON 4.41 1.1 3.43 1.1 3.43 0.56 3.59 0.56 3.59 0.16 3.71 0.16 3.71 0.62 3.49 0.62 3.49 1.04 4.17 1.04 4.17 0.485 4.18 0.485 4.18 0.425 4.24 0.425 4.24 0.545 4.23 0.545 4.23 1.04 4.41 1.04 ;
      POLYGON 4.04 0.94 3.59 0.94 3.59 0.88 3.98 0.88 3.98 0.4 4.04 0.4 ;
      POLYGON 3.945 1.26 3.27 1.26 3.27 0.23 3.03 0.23 3.03 0.17 3.33 0.17 3.33 1.2 3.945 1.2 ;
      RECT 3.09 0.695 3.17 1.195 ;
      POLYGON 2.77 0.495 2.69 0.495 2.69 0.25 2.515 0.25 2.515 0.17 2.77 0.17 ;
      POLYGON 2.59 1.245 2.305 1.245 2.305 1.315 2.245 1.315 2.245 1.245 1.465 1.245 1.465 1.185 2.53 1.185 2.53 0.465 2.47 0.465 2.47 0.405 2.59 0.405 ;
      POLYGON 2.27 0.805 1.895 0.805 1.895 0.56 1.975 0.56 1.975 0.725 2.27 0.725 ;
      POLYGON 1.8 1.025 1.365 1.025 1.365 1.15 0.34 1.15 0.34 0.73 0.4 0.73 0.4 1.09 1.305 1.09 1.305 0.965 1.735 0.965 1.735 0.465 1.675 0.465 1.675 0.405 1.795 0.405 1.795 0.905 1.8 0.905 ;
      POLYGON 0.56 0.78 0.5 0.78 0.5 0.63 0.165 0.63 0.165 1.29 0.105 1.29 0.105 0.57 0.18 0.57 0.18 0.49 0.31 0.49 0.31 0.57 0.56 0.57 ;
  END
END DLY4X4

MACRO EDFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFHQX1 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.603775 LAYER Metal1 ;
    ANTENNADIFFAREA 3.01475 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2601 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.010669 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 79.48673575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.18 1.09 3.06 1.09 3.06 0.79 3.1 0.79 3.1 0.535 3.18 0.535 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.5643565 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.765 0.715 4.555 0.715 4.555 0.685 4.245 0.685 4.245 0.745 4.185 0.745 4.185 0.625 4.3 0.625 4.3 0.365 3.895 0.365 3.895 0.905 3.835 0.905 3.835 0.305 4.36 0.305 4.36 0.625 4.765 0.625 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.77 0.935 4.455 0.935 4.455 0.97 4.375 0.97 4.375 0.785 4.455 0.785 4.455 0.815 4.77 0.815 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.73 0.34 1.23 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 1.77 0 1.77 0 1.65 0.335 1.65 0.335 1.33 0.395 1.33 0.395 1.65 1.68 1.65 1.68 1.19 1.74 1.19 1.74 1.65 2.825 1.65 2.825 1.35 2.945 1.35 2.945 1.41 2.885 1.41 2.885 1.65 3.495 1.65 3.495 1.35 3.615 1.35 3.615 1.41 3.555 1.41 3.555 1.65 4.43 1.65 4.43 1.245 4.49 1.245 4.49 1.65 5 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 0.06 4.52 0.06 4.52 0.525 4.46 0.525 4.46 0.06 3.5 0.06 3.5 0.49 3.44 0.49 3.44 0.06 2.78 0.06 2.78 0.425 2.84 0.425 2.84 0.485 2.72 0.485 2.72 0.06 1.74 0.06 1.74 0.19 1.8 0.19 1.8 0.25 1.68 0.25 1.68 0.06 0.435 0.06 0.435 0.465 0.375 0.465 0.375 0.06 0 0.06 0 -0.06 5 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.93 1.13 4.725 1.13 4.725 1.19 4.665 1.19 4.665 1.13 4.215 1.13 4.215 0.905 4.155 0.905 4.155 0.845 4.275 0.845 4.275 1.07 4.87 1.07 4.87 0.525 4.665 0.525 4.665 0.405 4.725 0.405 4.725 0.465 4.93 0.465 ;
      POLYGON 4.2 0.525 4.055 0.525 4.055 1.365 3.995 1.365 3.995 1.25 2.68 1.25 2.68 1.28 1.9 1.28 1.9 1.09 1.58 1.09 1.58 1.28 1.045 1.28 1.045 1.06 0.87 1.06 0.87 0.57 0.81 0.57 0.81 0.51 0.93 0.51 0.93 1 1.105 1 1.105 1.22 1.52 1.22 1.52 1.03 1.96 1.03 1.96 1.22 2.62 1.22 2.62 1.19 3.995 1.19 3.995 0.465 4.2 0.465 ;
      POLYGON 3.88 1.065 3.675 1.065 3.675 0.865 3.28 0.865 3.28 0.805 3.675 0.805 3.675 0.545 3.615 0.545 3.615 0.485 3.735 0.485 3.735 1.005 3.88 1.005 ;
      POLYGON 3.575 0.705 3.28 0.705 3.28 0.435 3 0.435 3 0.645 2.745 0.645 2.745 1.06 2.52 1.06 2.52 1.12 2.46 1.12 2.46 1 2.685 1 2.685 0.645 2.44 0.645 2.44 0.48 2.5 0.48 2.5 0.585 2.94 0.585 2.94 0.375 3.34 0.375 3.34 0.645 3.575 0.645 ;
      POLYGON 2.585 0.9 2.525 0.9 2.525 0.805 2.295 0.805 2.295 0.79 2.22 0.79 2.22 0.73 2.28 0.73 2.28 0.41 1.47 0.41 1.47 0.77 1.41 0.77 1.41 0.41 1.09 0.41 1.09 0.84 1.15 0.84 1.15 0.9 1.03 0.9 1.03 0.41 0.7 0.41 0.7 0.79 0.6 0.79 0.6 1.355 0.54 1.355 0.54 0.73 0.64 0.73 0.64 0.35 2.34 0.35 2.34 0.745 2.585 0.745 ;
      POLYGON 2.18 0.57 2.12 0.57 2.12 1.12 2.06 1.12 2.06 0.93 1.73 0.93 1.73 0.81 1.79 0.81 1.79 0.87 2.06 0.87 2.06 0.51 2.18 0.51 ;
      POLYGON 1.96 0.77 1.9 0.77 1.9 0.71 1.63 0.71 1.63 0.93 1.31 0.93 1.31 1.12 1.25 1.12 1.25 0.57 1.19 0.57 1.19 0.51 1.31 0.51 1.31 0.87 1.57 0.87 1.57 0.65 1.96 0.65 ;
      POLYGON 0.54 0.63 0.16 0.63 0.16 1.31 0.19 1.31 0.19 1.43 0.13 1.43 0.13 1.37 0.1 1.37 0.1 0.57 0.17 0.57 0.17 0.37 0.23 0.37 0.23 0.57 0.54 0.57 ;
  END
END EDFFHQX1

MACRO EDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFHQX2 0 0 ;
  SIZE 5.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.76715 LAYER Metal1 ;
    ANTENNADIFFAREA 3.42475 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.295425 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.36667525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 73.22670725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.175 1.14 3.045 1.14 3.045 0.92 2.86 0.92 2.86 0.79 3.045 0.79 3.045 0.55 3.165 0.55 3.165 0.63 3.125 0.63 3.125 1.06 3.175 1.06 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 16.5346535 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.94 0.73 4.86 0.73 4.86 0.66 4.17 0.66 4.17 0.8 4.11 0.8 4.11 0.6 4.235 0.6 4.235 0.34 3.85 0.34 3.85 0.98 3.79 0.98 3.79 0.28 4.295 0.28 4.295 0.6 4.94 0.6 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.76 0.84 4.54 0.84 4.54 1.03 4.46 1.03 4.46 0.84 4.45 0.84 4.45 0.76 4.76 0.76 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.425 1.13 0.235 1.13 0.235 1.085 0.23 1.085 0.23 0.745 0.31 0.745 0.31 1.005 0.425 1.005 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.2 1.77 0 1.77 0 1.65 0.295 1.65 0.295 1.23 0.355 1.23 0.355 1.65 1.685 1.65 1.685 1.3 1.625 1.3 1.625 1.24 1.745 1.24 1.745 1.65 2.82 1.65 2.82 1.4 2.94 1.4 2.94 1.46 2.88 1.46 2.88 1.65 3.29 1.65 3.29 1.4 3.41 1.4 3.41 1.46 3.35 1.46 3.35 1.65 4.535 1.65 4.535 1.29 4.595 1.29 4.595 1.65 5.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.2 0.06 4.595 0.06 4.595 0.5 4.535 0.5 4.535 0.06 3.485 0.06 3.485 0.5 3.425 0.5 3.425 0.06 2.785 0.06 2.785 0.5 2.725 0.5 2.725 0.06 1.685 0.06 1.685 0.41 1.745 0.41 1.745 0.47 1.625 0.47 1.625 0.06 0.325 0.06 0.325 0.4 0.385 0.4 0.385 0.46 0.265 0.46 0.265 0.06 0 0.06 0 -0.06 5.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.1 1.19 4.995 1.19 4.995 1.315 4.935 1.315 4.935 1.19 4.29 1.19 4.29 0.86 4.35 0.86 4.35 1.13 5.04 1.13 5.04 0.5 4.935 0.5 4.935 0.38 4.995 0.38 4.995 0.44 5.1 0.44 ;
      POLYGON 4.135 0.5 4.01 0.5 4.01 1.41 3.95 1.41 3.95 1.3 1.845 1.3 1.845 1.14 1.525 1.14 1.525 1.3 0.92 1.3 0.92 1.08 0.745 1.08 0.745 0.555 0.685 0.555 0.685 0.495 0.805 0.495 0.805 1.02 0.98 1.02 0.98 1.24 1.465 1.24 1.465 1.08 1.905 1.08 1.905 1.24 3.95 1.24 3.95 0.44 4.135 0.44 ;
      POLYGON 3.75 1.14 3.63 1.14 3.63 0.96 3.225 0.96 3.225 0.84 3.285 0.84 3.285 0.9 3.63 0.9 3.63 0.52 3.69 0.52 3.69 1.08 3.75 1.08 ;
      POLYGON 3.53 0.8 3.47 0.8 3.47 0.74 3.265 0.74 3.265 0.45 2.945 0.45 2.945 0.66 2.7 0.66 2.7 1.08 2.475 1.08 2.475 1.14 2.415 1.14 2.415 1.02 2.64 1.02 2.64 0.66 2.385 0.66 2.385 0.465 2.445 0.465 2.445 0.6 2.885 0.6 2.885 0.39 3.325 0.39 3.325 0.68 3.53 0.68 ;
      POLYGON 2.54 0.92 2.48 0.92 2.48 0.86 2.225 0.86 2.225 0.715 2.165 0.715 2.165 0.655 2.225 0.655 2.225 0.395 1.905 0.395 1.905 0.63 1.465 0.63 1.465 0.395 1.345 0.395 1.345 0.755 1.285 0.755 1.285 0.395 0.965 0.395 0.965 0.86 1.025 0.86 1.025 0.92 0.905 0.92 0.905 0.395 0.585 0.395 0.585 1.255 0.525 1.255 0.525 0.525 0.515 0.525 0.515 0.335 1.525 0.335 1.525 0.57 1.845 0.57 1.845 0.335 2.285 0.335 2.285 0.8 2.54 0.8 ;
      POLYGON 2.125 0.555 2.065 0.555 2.065 1.14 2.005 1.14 2.005 0.95 1.605 0.95 1.605 0.89 2.005 0.89 2.005 0.495 2.125 0.495 ;
      POLYGON 1.905 0.79 1.505 0.79 1.505 0.915 1.185 0.915 1.185 1.14 1.125 1.14 1.125 0.555 1.065 0.555 1.065 0.495 1.185 0.495 1.185 0.855 1.445 0.855 1.445 0.73 1.905 0.73 ;
      POLYGON 0.425 0.645 0.13 0.645 0.13 1.255 0.07 1.255 0.07 0.395 0.13 0.395 0.13 0.585 0.425 0.585 ;
  END
END EDFFHQX2

MACRO EDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFHQX4 0 0 ;
  SIZE 6.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.320775 LAYER Metal1 ;
    ANTENNADIFFAREA 4.0591 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.371025 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.950273 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 70.27289275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.9 0.63 3.84 0.63 3.84 0.81 3.14 0.81 3.14 1.005 3.225 1.005 3.225 1.125 3.725 1.125 3.725 1.185 3.17 1.185 3.17 1.16 3.165 1.16 3.165 1.085 3.035 1.085 3.035 1.005 3.08 1.005 3.08 0.63 3.02 0.63 3.02 0.57 3.14 0.57 3.14 0.75 3.78 0.75 3.78 0.57 3.9 0.57 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 15.280528 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.965 0.705 5.835 0.705 5.835 0.545 5.36 0.545 5.36 0.685 5.24 0.685 5.24 0.625 5.3 0.625 5.3 0.305 4.98 0.305 4.98 0.915 4.92 0.915 4.92 0.245 5.36 0.245 5.36 0.485 5.895 0.485 5.895 0.625 5.965 0.625 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.735 0.95 5.46 0.95 5.46 0.79 5.655 0.79 5.655 0.645 5.735 0.645 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.81 0.34 1.31 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 0 1.77 0 1.65 0.365 1.65 0.365 1.51 0.425 1.51 0.425 1.65 1.75 1.65 1.75 1.23 1.81 1.23 1.81 1.65 2.9 1.65 2.9 1.445 3.02 1.445 3.02 1.505 2.96 1.505 2.96 1.65 3.37 1.65 3.37 1.445 3.49 1.445 3.49 1.505 3.43 1.505 3.43 1.65 3.87 1.65 3.87 1.51 3.93 1.51 3.93 1.65 4.355 1.65 4.355 1.51 4.415 1.51 4.415 1.65 5.515 1.65 5.515 1.225 5.575 1.225 5.575 1.65 6.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 5.575 0.06 5.575 0.385 5.515 0.385 5.515 0.06 4.66 0.06 4.66 0.2 4.6 0.2 4.6 0.06 4.22 0.06 4.22 0.52 4.16 0.52 4.16 0.06 3.52 0.06 3.52 0.49 3.4 0.49 3.4 0.43 3.46 0.43 3.46 0.06 2.76 0.06 2.76 0.555 2.7 0.555 2.7 0.06 1.75 0.06 1.75 0.27 1.63 0.27 1.63 0.21 1.69 0.21 1.69 0.06 0.45 0.06 0.45 0.55 0.39 0.55 0.39 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.125 1.11 5.97 1.11 5.97 1.17 5.91 1.17 5.91 1.11 5.3 1.11 5.3 0.885 5.24 0.885 5.24 0.825 5.36 0.825 5.36 1.05 6.065 1.05 6.065 0.525 5.995 0.525 5.995 0.405 6.055 0.405 6.055 0.465 6.125 0.465 ;
      POLYGON 5.2 0.525 5.14 0.525 5.14 1.345 1.91 1.345 1.91 1.13 1.65 1.13 1.65 1.32 0.995 1.32 0.995 1.1 0.82 1.1 0.82 0.55 0.94 0.55 0.94 0.61 0.88 0.61 0.88 1.04 1.055 1.04 1.055 1.26 1.59 1.26 1.59 1.07 1.97 1.07 1.97 1.285 5.08 1.285 5.08 0.465 5.14 0.465 5.14 0.405 5.2 0.405 ;
      POLYGON 4.935 1.135 4.875 1.135 4.875 1.075 4.48 1.075 4.48 1.025 4.18 1.025 4.18 1.16 4.12 1.16 4.12 1.025 3.54 1.025 3.54 0.91 3.66 0.91 3.66 0.965 4.48 0.965 4.48 0.525 4.365 0.525 4.365 0.405 4.425 0.405 4.425 0.465 4.76 0.465 4.76 0.405 4.82 0.405 4.82 0.525 4.54 0.525 4.54 1.015 4.935 1.015 ;
      POLYGON 4.38 0.77 4.145 0.77 4.145 0.865 4.025 0.865 4.025 0.805 4.085 0.805 4.085 0.705 4 0.705 4 0.47 3.68 0.47 3.68 0.65 3.24 0.65 3.24 0.47 2.92 0.47 2.92 0.715 2.715 0.715 2.715 1.135 2.39 1.135 2.39 1.075 2.655 1.075 2.655 0.715 2.39 0.715 2.39 0.52 2.45 0.52 2.45 0.655 2.86 0.655 2.86 0.41 3.3 0.41 3.3 0.59 3.62 0.59 3.62 0.41 4.06 0.41 4.06 0.645 4.145 0.645 4.145 0.71 4.38 0.71 ;
      POLYGON 2.555 0.975 2.495 0.975 2.495 0.875 2.23 0.875 2.23 0.43 1.48 0.43 1.48 0.81 1.395 0.81 1.395 0.69 1.42 0.69 1.42 0.43 1.1 0.43 1.1 0.94 1.04 0.94 1.04 0.43 0.72 0.43 0.72 0.89 0.66 0.89 0.66 1.385 0.6 1.385 0.6 0.83 0.66 0.83 0.66 0.55 0.595 0.55 0.595 0.37 2.29 0.37 2.29 0.815 2.555 0.815 ;
      POLYGON 2.13 1.185 2.07 1.185 2.07 0.97 1.74 0.97 1.74 0.85 1.8 0.85 1.8 0.91 2.07 0.91 2.07 0.59 2.01 0.59 2.01 0.53 2.13 0.53 ;
      POLYGON 1.97 0.81 1.91 0.81 1.91 0.75 1.64 0.75 1.64 0.97 1.26 0.97 1.26 1.16 1.2 1.16 1.2 0.53 1.32 0.53 1.32 0.59 1.26 0.59 1.26 0.91 1.58 0.91 1.58 0.69 1.97 0.69 ;
      POLYGON 0.56 0.73 0.44 0.73 0.44 0.71 0.16 0.71 0.16 1.48 0.1 1.48 0.1 0.65 0.185 0.65 0.185 0.455 0.245 0.455 0.245 0.65 0.56 0.65 ;
  END
END EDFFHQX4

MACRO EDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFHQX8 0 0 ;
  SIZE 6.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6975 LAYER Metal1 ;
    ANTENNADIFFAREA 4.5737 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.528525 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.99588475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 54.820491 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.5 0.66 3.14 0.66 3.14 0.965 4.345 0.965 4.345 1.025 2.995 1.025 2.995 0.965 3.06 0.965 3.06 0.79 3.08 0.79 3.08 0.66 3.03 0.66 3.03 0.54 3.09 0.54 3.09 0.6 3.5 0.6 3.5 0.54 3.56 0.54 3.56 0.6 3.97 0.6 3.97 0.54 4.03 0.54 4.03 0.6 4.44 0.6 4.44 0.54 4.5 0.54 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.30033 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.565 0.715 6.245 0.715 6.245 0.705 5.915 0.705 5.915 0.645 6.04 0.645 6.04 0.385 5.655 0.385 5.655 0.895 5.595 0.895 5.595 0.325 6.1 0.325 6.1 0.645 6.245 0.645 6.245 0.625 6.565 0.625 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.075 0.815 6.575 0.895 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.76 0.34 1.26 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.8 1.77 0 1.77 0 1.65 0.335 1.65 0.335 1.36 0.395 1.36 0.395 1.65 1.64 1.65 1.64 1.16 1.7 1.16 1.7 1.65 2.79 1.65 2.79 1.285 2.91 1.285 2.91 1.345 2.85 1.345 2.85 1.65 3.2 1.65 3.2 1.285 3.32 1.285 3.32 1.345 3.26 1.345 3.26 1.65 3.61 1.65 3.61 1.285 3.73 1.285 3.73 1.345 3.67 1.345 3.67 1.65 4.02 1.65 4.02 1.285 4.14 1.285 4.14 1.345 4.08 1.345 4.08 1.65 4.785 1.65 4.785 1.315 4.905 1.315 4.905 1.375 4.845 1.375 4.845 1.65 5.255 1.65 5.255 1.315 5.375 1.315 5.375 1.375 5.315 1.375 5.315 1.65 6.17 1.65 6.17 1.235 6.23 1.235 6.23 1.65 6.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.8 0.06 6.26 0.06 6.26 0.525 6.2 0.525 6.2 0.06 5.26 0.06 5.26 0.435 5.2 0.435 5.2 0.06 4.88 0.06 4.88 0.405 4.76 0.405 4.76 0.345 4.82 0.345 4.82 0.06 4.295 0.06 4.295 0.17 4.175 0.17 4.175 0.06 3.825 0.06 3.825 0.17 3.705 0.17 3.705 0.06 3.355 0.06 3.355 0.17 3.235 0.17 3.235 0.06 2.77 0.06 2.77 0.485 2.71 0.485 2.71 0.06 1.76 0.06 1.76 0.25 1.64 0.25 1.64 0.19 1.7 0.19 1.7 0.06 0.405 0.06 0.405 0.495 0.345 0.495 0.345 0.06 0 0.06 0 -0.06 6.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.735 1.055 6.465 1.055 6.465 1.115 6.405 1.115 6.405 1.055 5.915 1.055 5.915 0.805 5.975 0.805 5.975 0.995 6.675 0.995 6.675 0.525 6.405 0.525 6.405 0.405 6.465 0.405 6.465 0.465 6.735 0.465 ;
      POLYGON 5.94 0.545 5.815 0.545 5.815 1.355 5.755 1.355 5.755 1.215 4.24 1.215 4.24 1.185 2.69 1.185 2.69 1.25 1.8 1.25 1.8 1.06 1.54 1.06 1.54 1.25 1.005 1.25 1.005 1.03 0.83 1.03 0.83 0.54 0.77 0.54 0.77 0.48 0.89 0.48 0.89 0.97 1.065 0.97 1.065 1.19 1.48 1.19 1.48 1 1.86 1 1.86 1.19 2.63 1.19 2.63 1.125 4.3 1.125 4.3 1.155 5.755 1.155 5.755 0.485 5.94 0.485 ;
      POLYGON 5.61 1.055 4.995 1.055 4.995 0.865 3.98 0.865 3.98 0.8 4.1 0.8 4.1 0.805 4.995 0.805 4.995 0.455 5.055 0.455 5.055 0.535 5.375 0.535 5.375 0.485 5.495 0.485 5.495 0.545 5.435 0.545 5.435 0.595 5.055 0.595 5.055 0.995 5.61 0.995 ;
      POLYGON 4.895 0.705 4.6 0.705 4.6 0.44 2.93 0.44 2.93 0.645 2.725 0.645 2.725 1.025 2.53 1.025 2.53 1.06 2.41 1.06 2.41 1 2.47 1 2.47 0.965 2.665 0.965 2.665 0.645 2.4 0.645 2.4 0.45 2.46 0.45 2.46 0.585 2.87 0.585 2.87 0.38 4.66 0.38 4.66 0.645 4.895 0.645 ;
      POLYGON 2.565 0.865 2.505 0.865 2.505 0.805 2.26 0.805 2.26 0.795 2.23 0.795 2.23 0.675 2.24 0.675 2.24 0.38 1.92 0.38 1.92 0.41 1.43 0.41 1.43 0.74 1.37 0.74 1.37 0.38 1.05 0.38 1.05 0.64 1.11 0.64 1.11 0.87 1.05 0.87 1.05 0.7 0.99 0.7 0.99 0.38 0.67 0.38 0.67 1.325 0.6 1.325 0.6 1.385 0.54 1.385 0.54 1.265 0.61 1.265 0.61 0.495 0.55 0.495 0.55 0.32 1.43 0.32 1.43 0.35 1.86 0.35 1.86 0.32 2.3 0.32 2.3 0.745 2.565 0.745 ;
      POLYGON 2.14 0.54 2.08 0.54 2.08 1.09 2.02 1.09 2.02 0.9 1.69 0.9 1.69 0.78 1.75 0.78 1.75 0.84 2.02 0.84 2.02 0.48 2.14 0.48 ;
      POLYGON 1.92 0.74 1.86 0.74 1.86 0.68 1.59 0.68 1.59 0.9 1.27 0.9 1.27 1.09 1.21 1.09 1.21 0.54 1.15 0.54 1.15 0.48 1.27 0.48 1.27 0.84 1.53 0.84 1.53 0.62 1.92 0.62 ;
      POLYGON 0.51 0.66 0.16 0.66 0.16 1.36 0.19 1.36 0.19 1.48 0.13 1.48 0.13 1.42 0.1 1.42 0.1 0.6 0.14 0.6 0.14 0.4 0.2 0.4 0.2 0.6 0.51 0.6 ;
  END
END EDFFHQX8

MACRO EDFFTRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFTRX1 0 0 ;
  SIZE 7.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8841 LAYER Metal1 ;
    ANTENNADIFFAREA 4.00355 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.308475 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.591296 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 98.74544125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.01 0.64 1 0.64 1 1.16 0.94 1.16 0.94 0.73 0.86 0.73 0.86 0.6 0.95 0.6 0.95 0.505 1.01 0.505 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9342 LAYER Metal1 ;
    ANTENNADIFFAREA 4.00355 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.308475 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.75370775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 99.52832475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.325 1.29 0.245 1.29 0.245 0.73 0.06 0.73 0.06 0.6 0.245 0.6 0.245 0.54 0.325 0.54 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.94 1.11 6.735 1.11 6.735 0.98 6.86 0.98 6.86 0.735 6.94 0.735 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.365 0.895 6.235 0.895 6.235 0.87 5.83 0.87 5.83 0.79 6.365 0.79 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.94 1.14 4.86 1.14 4.86 0.87 4.71 0.87 4.71 0.79 4.94 0.79 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.35 1.06 1.34 1.06 1.34 1.19 1.26 1.19 1.26 0.98 1.27 0.98 1.27 0.7 1.35 0.7 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 1.77 0 1.77 0 1.65 0.5 1.65 0.5 1.285 0.56 1.285 0.56 1.65 1.155 1.65 1.155 1.45 1.275 1.45 1.275 1.51 1.215 1.51 1.215 1.65 1.965 1.65 1.965 1.185 2.01 1.185 2.01 1.125 2.07 1.125 2.07 1.245 2.025 1.245 2.025 1.65 3.015 1.65 3.015 1.51 3.075 1.51 3.075 1.65 3.91 1.65 3.91 1.49 4.03 1.49 4.03 1.55 3.97 1.55 3.97 1.65 4.835 1.65 4.835 1.51 4.895 1.51 4.895 1.65 6.785 1.65 6.785 1.37 6.845 1.37 6.845 1.65 7.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 0.06 6.815 0.06 6.815 0.635 6.755 0.635 6.755 0.06 5.76 0.06 5.76 0.31 5.82 0.31 5.82 0.37 5.7 0.37 5.7 0.06 5.505 0.06 5.505 0.31 5.565 0.31 5.565 0.37 5.445 0.37 5.445 0.06 5.05 0.06 5.05 0.37 4.93 0.37 4.93 0.31 4.99 0.31 4.99 0.06 4.11 0.06 4.11 0.17 3.99 0.17 3.99 0.06 3.13 0.06 3.13 0.375 3.19 0.375 3.19 0.435 3.07 0.435 3.07 0.06 2.11 0.06 2.11 0.545 1.99 0.545 1.99 0.485 2.05 0.485 2.05 0.06 1.215 0.06 1.215 0.6 1.155 0.6 1.155 0.06 0.56 0.06 0.56 0.2 0.5 0.2 0.5 0.06 0 0.06 0 -0.06 7.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.1 1.27 6.135 1.27 6.135 1.35 6 1.35 6 1.29 6.075 1.29 6.075 1.21 7.04 1.21 7.04 0.54 7.1 0.54 ;
      POLYGON 6.61 1.02 6.55 1.02 6.55 0.69 5.375 0.69 5.375 0.63 6.55 0.63 6.55 0.54 6.61 0.54 ;
      POLYGON 6.195 1.095 6.075 1.095 6.075 1.03 5.74 1.03 5.74 1.125 5.67 1.125 5.67 0.85 5.215 0.85 5.215 0.53 4.77 0.53 4.77 0.235 4.27 0.235 4.27 0.385 3.77 0.385 3.77 0.325 4.21 0.325 4.21 0.175 4.83 0.175 4.83 0.47 5.165 0.47 5.165 0.305 5.225 0.305 5.225 0.47 5.92 0.47 5.92 0.335 6.13 0.335 6.13 0.395 5.98 0.395 5.98 0.53 5.275 0.53 5.275 0.79 5.73 0.79 5.73 0.97 6.135 0.97 6.135 1.035 6.195 1.035 ;
      POLYGON 5.975 1.19 5.9 1.19 5.9 1.285 5.32 1.285 5.32 1.19 5.245 1.19 5.245 1.13 5.38 1.13 5.38 1.225 5.84 1.225 5.84 1.13 5.975 1.13 ;
      POLYGON 5.56 1.125 5.48 1.125 5.48 1.03 5.145 1.03 5.145 1.125 5.065 1.125 5.065 0.95 5.56 0.95 ;
      POLYGON 5.22 1.35 2.245 1.35 2.245 1.405 2.125 1.405 2.125 1.345 2.185 1.345 2.185 1.025 1.865 1.025 1.865 1.35 1.1 1.35 1.1 0.74 1.16 0.74 1.16 1.29 1.805 1.29 1.805 1.025 1.67 1.025 1.67 0.54 1.73 0.54 1.73 0.965 2.245 0.965 2.245 1.29 5.22 1.29 ;
      POLYGON 5.02 0.69 4.61 0.69 4.61 1.125 4.55 1.125 4.55 0.335 4.67 0.335 4.67 0.395 4.61 0.395 4.61 0.63 5.02 0.63 ;
      POLYGON 4.345 0.57 4.285 0.57 4.285 1.12 4.145 1.12 4.145 1.06 4.225 1.06 4.225 0.915 3.61 0.915 3.61 0.855 4.225 0.855 4.225 0.51 4.345 0.51 ;
      POLYGON 4.125 0.755 3.61 0.755 3.61 0.38 3.35 0.38 3.35 0.89 3.29 0.89 3.29 0.595 2.91 0.595 2.91 0.38 2.65 0.38 2.65 0.86 2.53 0.86 2.53 0.8 2.59 0.8 2.59 0.38 2.27 0.38 2.27 0.705 1.83 0.705 1.83 0.44 1.425 0.44 1.425 0.54 1.51 0.54 1.51 0.93 1.57 0.93 1.57 0.99 1.45 0.99 1.45 0.6 1.365 0.6 1.365 0.38 1.89 0.38 1.89 0.645 2.21 0.645 2.21 0.32 2.305 0.32 2.305 0.275 2.425 0.275 2.425 0.32 2.97 0.32 2.97 0.535 3.29 0.535 3.29 0.32 3.67 0.32 3.67 0.695 4.125 0.695 ;
      POLYGON 3.51 1.15 3.45 1.15 3.45 1.05 3.13 1.05 3.13 0.935 2.91 0.935 2.91 0.875 3.19 0.875 3.19 0.99 3.45 0.99 3.45 0.48 3.51 0.48 ;
      POLYGON 3.19 0.755 2.81 0.755 2.81 1.15 2.75 1.15 2.75 0.48 2.81 0.48 2.81 0.695 3.19 0.695 ;
      POLYGON 2.49 0.57 2.43 0.57 2.43 0.96 2.48 0.96 2.48 1.15 2.42 1.15 2.42 1.02 2.37 1.02 2.37 0.865 1.915 0.865 1.915 0.805 2.37 0.805 2.37 0.51 2.49 0.51 ;
      POLYGON 0.76 1.02 0.68 1.02 0.68 0.79 0.425 0.79 0.425 0.71 0.68 0.71 0.68 0.54 0.76 0.54 ;
  END
END EDFFTRX1

MACRO EDFFTRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFTRX2 0 0 ;
  SIZE 7.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.304125 LAYER Metal1 ;
    ANTENNADIFFAREA 4.5498 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.37305 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.5376625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 89.65822275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.215 1.11 7.06 1.11 7.06 0.98 7.065 0.98 7.065 0.54 7.145 0.54 7.145 1.03 7.215 1.03 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.304125 LAYER Metal1 ;
    ANTENNADIFFAREA 4.5498 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.37305 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.5376625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 89.65822275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.94 0.92 6.755 0.92 6.755 1.14 6.625 1.14 6.625 1.06 6.675 1.06 6.675 0.54 6.755 0.54 6.755 0.79 6.94 0.79 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.365 1.085 6.235 1.085 6.235 1.005 6.285 1.005 6.285 0.635 6.365 0.635 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.66 0.75 2.74 1.25 ;
    END
  END RN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.675926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.48 0.83 1.365 0.83 1.365 1.15 0.705 1.15 0.705 1.085 0.635 1.085 0.635 1.005 0.705 1.005 0.705 0.73 0.765 0.73 0.765 1.09 1.305 1.09 1.305 0.77 1.48 0.77 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 0.73 0.34 0.73 0.34 0.88 0.26 0.88 0.26 0.6 0.56 0.6 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.8 1.77 0 1.77 0 1.65 0.63 1.65 0.63 1.54 0.75 1.54 0.75 1.65 2.61 1.65 2.61 1.51 2.67 1.51 2.67 1.65 3.45 1.65 3.45 1.51 3.51 1.51 3.51 1.65 4.5 1.65 4.5 1.54 4.62 1.54 4.62 1.65 5.68 1.65 5.68 1.125 5.8 1.125 5.8 1.185 5.74 1.185 5.74 1.65 6.42 1.65 6.42 1.51 6.48 1.51 6.48 1.65 6.86 1.65 6.86 1.4 6.98 1.4 6.98 1.46 6.92 1.46 6.92 1.65 7.36 1.65 7.36 1.51 7.42 1.51 7.42 1.65 7.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.8 0.06 7.35 0.06 7.35 0.52 7.29 0.52 7.29 0.06 6.94 0.06 6.94 0.52 6.88 0.52 6.88 0.06 6.495 0.06 6.495 0.535 6.435 0.535 6.435 0.06 5.77 0.06 5.77 0.17 5.65 0.17 5.65 0.06 4.56 0.06 4.56 0.365 4.62 0.365 4.62 0.425 4.5 0.425 4.5 0.06 3.5 0.06 3.5 0.25 3.38 0.25 3.38 0.19 3.44 0.19 3.44 0.06 2.57 0.06 2.57 0.33 2.51 0.33 2.51 0.06 1.84 0.06 1.84 0.29 1.9 0.29 1.9 0.35 1.78 0.35 1.78 0.06 1.545 0.06 1.545 0.35 1.485 0.35 1.485 0.06 0.69 0.06 0.69 0.5 0.63 0.5 0.63 0.06 0 0.06 0 -0.06 7.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.585 1.12 7.525 1.12 7.525 0.815 7.245 0.815 7.245 0.755 7.525 0.755 7.525 0.54 7.585 0.54 ;
      POLYGON 7.58 1.385 7.52 1.385 7.52 1.325 7.08 1.325 7.08 1.3 5.975 1.3 5.975 1.36 5.905 1.36 5.905 1.025 5.58 1.025 5.58 1.41 2.39 1.41 2.39 1.47 2.33 1.47 2.33 1.35 5.52 1.35 5.52 0.965 5.905 0.965 5.905 0.57 6.025 0.57 6.025 0.63 5.965 0.63 5.965 1.24 6.465 1.24 6.465 0.9 6.515 0.9 6.515 0.7 6.575 0.7 6.575 0.96 6.525 0.96 6.525 1.24 7.14 1.24 7.14 1.265 7.58 1.265 ;
      POLYGON 6.29 0.535 6.185 0.535 6.185 0.905 6.135 0.905 6.135 1.12 6.075 1.12 6.075 0.845 6.125 0.845 6.125 0.47 5.49 0.47 5.49 0.385 5.1 0.385 5.1 0.905 4.98 0.905 4.98 0.845 5.04 0.845 5.04 0.385 4.78 0.385 4.78 0.585 4.315 0.585 4.315 0.85 4.255 0.85 4.255 0.415 3.88 0.415 3.88 0.76 3.395 0.76 3.395 0.7 3.82 0.7 3.82 0.355 4.315 0.355 4.315 0.525 4.72 0.525 4.72 0.325 5.355 0.325 5.355 0.16 5.475 0.16 5.475 0.325 5.55 0.325 5.55 0.41 6.29 0.41 ;
      POLYGON 5.805 0.845 5.745 0.845 5.745 0.705 5.26 0.705 5.26 1.09 5.14 1.09 5.14 1.03 5.2 1.03 5.2 0.645 5.33 0.645 5.33 0.485 5.39 0.485 5.39 0.645 5.805 0.645 ;
      POLYGON 5.48 0.865 5.42 0.865 5.42 1.25 3.935 1.25 3.935 0.93 3.345 0.93 3.345 1.12 3.285 1.12 3.285 0.93 3.235 0.93 3.235 0.575 3 0.575 3 0.515 3.295 0.515 3.295 0.87 3.995 0.87 3.995 1.19 5.36 1.19 5.36 0.805 5.48 0.805 ;
      POLYGON 4.94 0.745 4.88 0.745 4.88 1.03 4.94 1.03 4.94 1.09 4.82 1.09 4.82 0.745 4.415 0.745 4.415 0.685 4.88 0.685 4.88 0.485 4.94 0.485 ;
      POLYGON 4.715 0.93 4.655 0.93 4.655 1.01 4.215 1.01 4.215 1.09 4.095 1.09 4.095 0.575 3.98 0.575 3.98 0.515 4.155 0.515 4.155 0.95 4.595 0.95 4.595 0.87 4.715 0.87 ;
      POLYGON 3.72 0.39 3.66 0.39 3.66 0.41 3.22 0.41 3.22 0.295 2.73 0.295 2.73 0.49 2.335 0.49 2.335 0.67 1.76 0.67 1.76 1.02 1.7 1.02 1.7 0.67 1.205 0.67 1.205 0.99 1.085 0.99 1.085 0.93 1.145 0.93 1.145 0.54 1.205 0.54 1.205 0.61 2.275 0.61 2.275 0.37 2.335 0.37 2.335 0.43 2.67 0.43 2.67 0.235 3.28 0.235 3.28 0.35 3.6 0.35 3.6 0.33 3.72 0.33 ;
      POLYGON 2.9 1.03 2.84 1.03 2.84 0.65 2.51 0.65 2.51 0.71 2.45 0.71 2.45 0.59 2.83 0.59 2.83 0.395 2.89 0.395 2.89 0.59 2.9 0.59 ;
      POLYGON 2.435 1.03 2.355 1.03 2.355 0.905 2.045 0.905 2.045 1.03 1.965 1.03 1.965 0.825 2.435 0.825 ;
      POLYGON 2.23 1.19 1.525 1.19 1.525 1.085 1.465 1.085 1.465 1.025 1.585 1.025 1.585 1.13 2.17 1.13 2.17 1.005 2.23 1.005 ;
      POLYGON 2.12 0.3 2.06 0.3 2.06 0.51 1.325 0.51 1.325 0.44 0.925 0.44 0.925 0.93 0.985 0.93 0.985 0.99 0.865 0.99 0.865 0.38 1.385 0.38 1.385 0.45 2 0.45 2 0.24 2.12 0.24 ;
      POLYGON 1.31 1.31 0.425 1.31 0.425 1.04 0.1 1.04 0.1 0.44 0.425 0.44 0.425 0.38 0.485 0.38 0.485 0.5 0.16 0.5 0.16 0.98 0.485 0.98 0.485 1.25 1.31 1.25 ;
  END
END EDFFTRX2

MACRO EDFFTRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFTRX4 0 0 ;
  SIZE 8.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6578 LAYER Metal1 ;
    ANTENNADIFFAREA 5.1215 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.5202 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.953864 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 70.35755475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.89 0.99 7.28 0.99 7.28 0.92 7.26 0.92 7.26 0.79 7.28 0.79 7.28 0.435 7.345 0.435 7.345 0.515 7.695 0.515 7.695 0.435 7.755 0.435 7.755 0.575 7.34 0.575 7.34 0.93 7.89 0.93 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6578 LAYER Metal1 ;
    ANTENNADIFFAREA 5.1215 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.5202 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.953864 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 70.35755475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.95 0.99 6.36 0.99 6.36 0.93 6.66 0.93 6.66 0.575 6.465 0.575 6.465 0.435 6.525 0.435 6.525 0.515 6.875 0.515 6.875 0.435 6.935 0.435 6.935 0.575 6.72 0.575 6.72 0.79 6.74 0.79 6.74 0.93 6.95 0.93 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.66 0.96 5.41 0.96 5.41 0.88 5.435 0.88 5.435 0.63 5.655 0.63 5.655 0.815 5.66 0.815 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.11 0.895 2.965 0.895 2.965 0.965 2.68 0.965 2.68 0.815 3.11 0.815 ;
    END
  END RN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 15.18518525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.45 0.92 1.365 0.92 1.365 1.275 0.635 1.275 0.635 1.195 0.705 1.195 0.705 0.805 0.765 0.805 0.765 1.215 1.305 1.215 1.305 0.86 1.45 0.86 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.605 0.92 0.34 0.92 0.34 0.97 0.26 0.97 0.26 0.79 0.525 0.79 0.525 0.735 0.605 0.735 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.4 1.77 0 1.77 0 1.65 0.63 1.65 0.63 1.54 0.75 1.54 0.75 1.65 2.545 1.65 2.545 1.51 2.605 1.51 2.605 1.65 2.94 1.65 2.94 1.51 3 1.51 3 1.65 3.805 1.65 3.805 1.51 3.865 1.51 3.865 1.65 4.825 1.65 4.825 1.54 4.945 1.54 4.945 1.65 5.725 1.65 5.725 1.54 5.845 1.54 5.845 1.65 6.125 1.65 6.125 1.25 6.245 1.25 6.245 1.31 6.185 1.31 6.185 1.65 6.595 1.65 6.595 1.25 6.715 1.25 6.715 1.31 6.655 1.31 6.655 1.65 7.065 1.65 7.065 1.25 7.185 1.25 7.185 1.31 7.125 1.31 7.125 1.65 7.535 1.65 7.535 1.25 7.655 1.25 7.655 1.31 7.595 1.31 7.595 1.65 8.005 1.65 8.005 1.25 8.125 1.25 8.125 1.31 8.065 1.31 8.065 1.65 8.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.4 0.06 7.965 0.06 7.965 0.415 7.905 0.415 7.905 0.06 7.55 0.06 7.55 0.415 7.49 0.415 7.49 0.06 7.14 0.06 7.14 0.415 7.08 0.415 7.08 0.06 6.73 0.06 6.73 0.415 6.67 0.415 6.67 0.06 6.32 0.06 6.32 0.415 6.26 0.415 6.26 0.06 5.83 0.06 5.83 0.47 5.77 0.47 5.77 0.06 4.77 0.06 4.77 0.545 4.83 0.545 4.83 0.605 4.71 0.605 4.71 0.06 3.75 0.06 3.75 0.39 3.81 0.39 3.81 0.45 3.69 0.45 3.69 0.06 2.815 0.06 2.815 0.17 2.695 0.17 2.695 0.06 2.35 0.06 2.35 0.2 2.29 0.2 2.29 0.06 1.69 0.06 1.69 0.38 1.75 0.38 1.75 0.44 1.63 0.44 1.63 0.06 1.53 0.06 1.53 0.44 1.41 0.44 1.41 0.38 1.47 0.38 1.47 0.06 0.69 0.06 0.69 0.635 0.63 0.635 0.63 0.06 0 0.06 0 -0.06 8.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 8.33 1.29 8.27 1.29 8.27 0.605 7.915 0.605 7.915 0.725 7.855 0.725 7.855 0.545 8.11 0.545 8.11 0.435 8.17 0.435 8.17 0.545 8.33 0.545 ;
      POLYGON 8.095 1.15 5.98 1.15 5.98 1.28 5.93 1.28 5.93 1.44 4.745 1.44 4.745 1.43 4.23 1.43 4.23 1.305 2.325 1.305 2.325 1.365 2.265 1.365 2.265 1.245 4.29 1.245 4.29 1.37 4.785 1.37 4.785 1.38 5.87 1.38 5.87 1.22 5.92 1.22 5.92 0.9 6.005 0.9 6.005 0.435 6.065 0.435 6.065 0.675 6.415 0.675 6.415 0.735 6.065 0.735 6.065 0.96 5.98 0.96 5.98 1.09 8.035 1.09 8.035 0.705 8.095 0.705 ;
      POLYGON 5.905 0.8 5.82 0.8 5.82 1.12 5.77 1.12 5.77 1.28 4.845 1.28 4.845 1.27 4.39 1.27 4.39 0.54 4.45 0.54 4.45 1.21 4.885 1.21 4.885 1.22 5.71 1.22 5.71 1.06 5.76 1.06 5.76 0.74 5.845 0.74 5.845 0.68 5.905 0.68 ;
      POLYGON 5.61 1.12 5.25 1.12 5.25 0.47 5.52 0.47 5.52 0.37 4.99 0.37 4.99 0.765 4.55 0.765 4.55 0.44 4.29 0.44 4.29 0.95 4.23 0.95 4.23 0.44 3.97 0.44 3.97 0.61 3.43 0.61 3.43 0.95 3.37 0.95 3.37 0.435 3.255 0.435 3.255 0.375 3.43 0.375 3.43 0.55 3.91 0.55 3.91 0.38 4.475 0.38 4.475 0.205 4.595 0.205 4.595 0.38 4.61 0.38 4.61 0.705 4.93 0.705 4.93 0.435 4.87 0.435 4.87 0.31 5.58 0.31 5.58 0.53 5.31 0.53 5.31 1.06 5.61 1.06 ;
      POLYGON 5.15 1.09 5 1.09 5 1.03 5.09 1.03 5.09 0.93 4.55 0.93 4.55 0.87 5.09 0.87 5.09 0.54 5.15 0.54 ;
      POLYGON 4.13 1.12 4.07 1.12 4.07 0.99 3.75 0.99 3.75 0.93 3.69 0.93 3.69 0.87 3.81 0.87 3.81 0.93 4.07 0.93 4.07 0.54 4.13 0.54 ;
      POLYGON 3.97 0.83 3.91 0.83 3.91 0.77 3.59 0.77 3.59 1.11 3.21 1.11 3.21 0.63 3.15 0.63 3.15 0.57 3.27 0.57 3.27 1.05 3.53 1.05 3.53 0.71 3.97 0.71 ;
      POLYGON 3.035 0.435 2.185 0.435 2.185 0.76 1.76 0.76 1.76 1.11 1.7 1.11 1.7 0.76 1.15 0.76 1.15 1.02 1.205 1.02 1.205 1.08 1.085 1.08 1.085 1.02 1.09 1.02 1.09 0.63 1.03 0.63 1.03 0.57 1.15 0.57 1.15 0.7 2.125 0.7 2.125 0.375 3.035 0.375 ;
      POLYGON 2.795 1.125 2.52 1.125 2.52 0.805 2.42 0.805 2.42 0.745 2.52 0.745 2.52 0.63 2.46 0.63 2.46 0.57 2.58 0.57 2.58 1.065 2.795 1.065 ;
      POLYGON 2.37 1.11 2.29 1.11 2.29 0.985 1.98 0.985 1.98 1.11 1.9 1.11 1.9 0.905 2.37 0.905 ;
      POLYGON 2.165 1.27 1.525 1.27 1.525 1.175 1.465 1.175 1.465 1.115 1.585 1.115 1.585 1.21 2.105 1.21 2.105 1.085 2.165 1.085 ;
      POLYGON 1.97 0.435 1.91 0.435 1.91 0.6 1.25 0.6 1.25 0.47 0.895 0.47 0.895 0.575 0.925 0.575 0.925 1.005 0.985 1.005 0.985 1.065 0.865 1.065 0.865 0.635 0.835 0.635 0.835 0.41 1.31 0.41 1.31 0.54 1.85 0.54 1.85 0.375 1.97 0.375 ;
      POLYGON 1.28 1.435 0.425 1.435 0.425 1.13 0.1 1.13 0.1 0.575 0.425 0.575 0.425 0.515 0.485 0.515 0.485 0.635 0.16 0.635 0.16 1.07 0.485 1.07 0.485 1.375 1.28 1.375 ;
  END
END EDFFTRX4

MACRO EDFFTRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFTRXL 0 0 ;
  SIZE 6.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5986 LAYER Metal1 ;
    ANTENNADIFFAREA 3.69445 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2754 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.066812 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 101.6122005 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.52 0.94 1.02 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6386 LAYER Metal1 ;
    ANTENNADIFFAREA 3.69445 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2754 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.21205525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 102.24400875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.285 1.02 0.205 1.02 0.205 0.73 0.06 0.73 0.06 0.6 0.205 0.6 0.205 0.54 0.285 0.54 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.435 1.11 6.26 1.11 6.26 0.855 6.23 0.855 6.23 0.735 6.435 0.735 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.388889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.965 0.895 5.835 0.895 5.835 0.845 5.405 0.845 5.405 0.765 5.965 0.765 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.54 1.18 4.46 1.18 4.46 0.93 4.29 0.93 4.29 0.85 4.54 0.85 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.165 1.02 1.085 1.02 1.085 0.77 1.06 0.77 1.06 0.545 1.14 0.545 1.14 0.69 1.165 0.69 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.8 1.77 0 1.77 0 1.65 0.495 1.65 0.495 1.285 0.555 1.285 0.555 1.65 1.115 1.65 1.115 1.295 1.175 1.295 1.175 1.65 1.64 1.65 1.64 1.155 1.725 1.155 1.725 1.095 1.785 1.095 1.785 1.215 1.7 1.215 1.7 1.65 2.65 1.65 2.65 1.49 2.77 1.49 2.77 1.55 2.71 1.55 2.71 1.65 3.54 1.65 3.54 1.49 3.66 1.49 3.66 1.55 3.6 1.55 3.6 1.65 4.415 1.65 4.415 1.51 4.475 1.51 4.475 1.65 6.3 1.65 6.3 1.37 6.36 1.37 6.36 1.65 6.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.8 0.06 6.33 0.06 6.33 0.635 6.27 0.635 6.27 0.06 5.39 0.06 5.39 0.285 5.45 0.285 5.45 0.345 5.33 0.345 5.33 0.06 5.115 0.06 5.115 0.285 5.175 0.285 5.175 0.345 5.055 0.345 5.055 0.06 4.63 0.06 4.63 0.43 4.51 0.43 4.51 0.37 4.57 0.37 4.57 0.06 3.715 0.06 3.715 0.17 3.595 0.17 3.595 0.06 2.775 0.06 2.775 0.42 2.835 0.42 2.835 0.48 2.715 0.48 2.715 0.06 1.84 0.06 1.84 0.2 1.78 0.2 1.78 0.06 1.155 0.06 1.155 0.2 1.095 0.2 1.095 0.06 0.555 0.06 0.555 0.2 0.495 0.2 0.495 0.06 0 0.06 0 -0.06 6.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.595 1.27 5.93 1.27 5.93 1.325 5.575 1.325 5.575 1.265 5.87 1.265 5.87 1.21 6.535 1.21 6.535 0.54 6.595 0.54 ;
      POLYGON 6.125 1.02 6.065 1.02 6.065 0.665 4.95 0.665 4.95 0.605 6.065 0.605 6.065 0.54 6.125 0.54 ;
      POLYGON 5.77 1.07 5.65 1.07 5.65 1.005 5.315 1.005 5.315 1.1 5.245 1.1 5.245 0.825 4.79 0.825 4.79 0.59 4.35 0.59 4.35 0.295 4.03 0.295 4.03 0.445 3.425 0.445 3.425 0.385 3.97 0.385 3.97 0.235 4.41 0.235 4.41 0.53 4.745 0.53 4.745 0.365 4.805 0.365 4.805 0.445 5.55 0.445 5.55 0.34 5.67 0.34 5.67 0.28 5.73 0.28 5.73 0.4 5.61 0.4 5.61 0.505 4.85 0.505 4.85 0.765 5.305 0.765 5.305 0.945 5.71 0.945 5.71 1.01 5.77 1.01 ;
      POLYGON 5.55 1.165 5.475 1.165 5.475 1.26 4.895 1.26 4.895 1.165 4.82 1.165 4.82 1.105 4.955 1.105 4.955 1.2 5.415 1.2 5.415 1.105 5.55 1.105 ;
      POLYGON 5.135 1.1 5.055 1.1 5.055 1.005 4.72 1.005 4.72 1.1 4.64 1.1 4.64 0.925 5.135 0.925 ;
      POLYGON 4.795 1.34 1.945 1.34 1.945 1.375 1.8 1.375 1.8 1.315 1.885 1.315 1.885 0.995 1.54 0.995 1.54 1.18 1.015 1.18 1.015 1.245 0.895 1.245 0.895 1.185 0.955 1.185 0.955 1.12 1.46 1.12 1.46 0.54 1.52 0.54 1.52 0.935 1.945 0.935 1.945 1.28 4.795 1.28 ;
      POLYGON 4.67 0.75 4.19 0.75 4.19 1.1 4.13 1.1 4.13 0.395 4.25 0.395 4.25 0.455 4.19 0.455 4.19 0.69 4.67 0.69 ;
      POLYGON 3.915 1.12 3.775 1.12 3.775 1.06 3.855 1.06 3.855 0.95 3.265 0.95 3.265 0.89 3.855 0.89 3.855 0.63 3.775 0.63 3.775 0.57 3.915 0.57 ;
      POLYGON 3.755 0.79 3.265 0.79 3.265 0.44 3.005 0.44 3.005 0.96 2.945 0.96 2.945 0.64 2.555 0.64 2.555 0.44 2.295 0.44 2.295 0.95 2.235 0.95 2.235 0.44 1.32 0.44 1.32 0.6 1.325 0.6 1.325 1.02 1.265 1.02 1.265 0.635 1.26 0.635 1.26 0.38 1.94 0.38 1.94 0.265 2.06 0.265 2.06 0.38 2.615 0.38 2.615 0.58 2.945 0.58 2.945 0.38 3.325 0.38 3.325 0.73 3.755 0.73 ;
      POLYGON 3.165 1.18 3.105 1.18 3.105 1.12 2.785 1.12 2.785 0.96 2.555 0.96 2.555 0.9 2.845 0.9 2.845 1.06 3.105 1.06 3.105 0.54 3.165 0.54 ;
      POLYGON 2.845 0.8 2.455 0.8 2.455 1.12 2.335 1.12 2.335 1.06 2.395 1.06 2.395 0.54 2.455 0.54 2.455 0.74 2.845 0.74 ;
      POLYGON 2.135 1.15 2.075 1.15 2.075 0.8 1.62 0.8 1.62 0.74 2.075 0.74 2.075 0.63 2.015 0.63 2.015 0.57 2.135 0.57 ;
      POLYGON 0.72 1.02 0.64 1.02 0.64 0.81 0.385 0.81 0.385 0.73 0.64 0.73 0.64 0.54 0.72 0.54 ;
  END
END EDFFTRXL

MACRO EDFFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFX1 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83885 LAYER Metal1 ;
    ANTENNADIFFAREA 3.2092 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.243675 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.65014875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 90.3170205 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.34 1.29 5.28 1.29 5.28 0.73 5.26 0.73 5.26 0.6 5.28 0.6 5.28 0.54 5.34 0.54 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.88645 LAYER Metal1 ;
    ANTENNADIFFAREA 3.2092 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.243675 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.845491 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 91.3388735 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.46 0.54 4.54 1.29 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 20 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.14 1.11 4.12 1.11 4.12 1.14 3.295 1.14 3.295 1.515 2.965 1.515 2.965 1.455 3.235 1.455 3.235 0.755 3.175 0.755 3.175 0.695 3.295 0.695 3.295 1.08 4.06 1.08 4.06 0.975 4.14 0.975 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.96 0.885 3.765 0.885 3.765 0.98 3.555 0.98 3.555 0.805 3.96 0.805 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 1.11 0.46 1.11 0.46 1.06 0.3 1.06 0.3 0.77 0.38 0.77 0.38 0.98 0.54 0.98 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 0 1.77 0 1.65 0.365 1.65 0.365 1.21 0.425 1.21 0.425 1.65 1.54 1.65 1.54 1.305 1.66 1.305 1.66 1.365 1.6 1.365 1.6 1.65 2.56 1.65 2.56 1.49 2.68 1.49 2.68 1.55 2.62 1.55 2.62 1.65 3.66 1.65 3.66 1.24 3.72 1.24 3.72 1.65 4.665 1.65 4.665 0.92 4.725 0.92 4.725 1.65 5.06 1.65 5.06 1.17 5.12 1.17 5.12 1.65 5.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5.105 0.06 5.105 0.2 5.045 0.2 5.045 0.06 4.86 0.06 4.86 0.2 4.8 0.2 4.8 0.06 3.72 0.06 3.72 0.19 3.78 0.19 3.78 0.25 3.66 0.25 3.66 0.06 2.68 0.06 2.68 0.575 2.62 0.575 2.62 0.06 1.66 0.06 1.66 0.22 1.54 0.22 1.54 0.16 1.6 0.16 1.6 0.06 0.425 0.06 0.425 0.51 0.365 0.51 0.365 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.125 0.795 4.98 0.795 4.98 1.02 4.9 1.02 4.9 0.54 4.98 0.54 4.98 0.715 5.125 0.715 ;
      POLYGON 4.7 0.82 4.64 0.82 4.64 0.385 3.94 0.385 3.94 0.41 2.915 0.41 2.915 1.01 2.855 1.01 2.855 1.11 2.915 1.11 2.915 1.17 2.795 1.17 2.795 1.01 2.58 1.01 2.58 0.89 2.64 0.89 2.64 0.95 2.855 0.95 2.855 0.35 3.88 0.35 3.88 0.325 4.7 0.325 ;
      POLYGON 4.3 1.27 4.28 1.27 4.28 1.33 4.22 1.33 4.22 1.21 4.24 1.21 4.24 0.705 3.455 0.705 3.455 0.89 3.395 0.89 3.395 0.645 4.24 0.645 4.24 0.545 4.105 0.545 4.105 0.485 4.3 0.485 ;
      POLYGON 3.255 0.57 3.075 0.57 3.075 1.21 3.12 1.21 3.12 1.33 1.76 1.33 1.76 1.205 1.44 1.205 1.44 1.33 1.015 1.33 1.015 1.205 0.84 1.205 0.84 0.54 0.9 0.54 0.9 1.145 1.075 1.145 1.075 1.27 1.38 1.27 1.38 1.145 1.82 1.145 1.82 1.27 3.015 1.27 3.015 0.51 3.255 0.51 ;
      POLYGON 2.755 0.79 2.48 0.79 2.48 1.16 2.155 1.16 2.155 1.1 2.42 1.1 2.42 0.78 2.24 0.78 2.24 0.54 2.3 0.54 2.3 0.72 2.755 0.72 ;
      POLYGON 2.32 1 2.26 1 2.26 0.94 2.08 0.94 2.08 0.855 1.995 0.855 1.995 0.735 2.08 0.735 2.08 0.415 1.06 0.415 1.06 0.86 1.12 0.86 1.12 0.92 1 0.92 1 0.415 0.7 0.415 0.7 1.235 0.64 1.235 0.64 0.355 1.26 0.355 1.26 0.295 1.38 0.295 1.38 0.355 2.14 0.355 2.14 0.88 2.32 0.88 ;
      POLYGON 1.98 0.635 1.895 0.635 1.895 0.955 1.98 0.955 1.98 1.17 1.92 1.17 1.92 1.015 1.445 1.015 1.445 0.92 1.565 0.92 1.565 0.955 1.835 0.955 1.835 0.575 1.92 0.575 1.92 0.515 1.98 0.515 ;
      POLYGON 1.735 0.8 1.28 0.8 1.28 1.17 1.22 1.17 1.22 0.63 1.16 0.63 1.16 0.57 1.28 0.57 1.28 0.74 1.735 0.74 ;
      POLYGON 0.54 0.73 0.48 0.73 0.48 0.67 0.2 0.67 0.2 1.235 0.14 1.235 0.14 0.415 0.2 0.415 0.2 0.61 0.54 0.61 ;
  END
END EDFFX1

MACRO EDFFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFX2 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.99235 LAYER Metal1 ;
    ANTENNADIFFAREA 3.284925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.30825 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.7075425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 74.97810225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.815 0.565 4.74 0.565 4.74 1.355 4.68 1.355 4.68 0.73 4.66 0.73 4.66 0.6 4.68 0.6 4.68 0.505 4.815 0.505 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.99235 LAYER Metal1 ;
    ANTENNADIFFAREA 3.284925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.30825 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.7075425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 74.97810225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.365 0.705 4.295 0.705 4.295 1.355 4.235 1.355 4.235 0.565 4.225 0.565 4.225 0.505 4.345 0.505 4.345 0.625 4.365 0.625 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 24.074074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.965 0.895 3.92 0.895 3.92 1.31 2.865 1.31 2.865 1.485 2.745 1.485 2.745 1.425 2.805 1.425 2.805 1.25 3.015 1.25 3.015 0.725 2.955 0.725 2.955 0.665 3.075 0.665 3.075 1.25 3.86 1.25 3.86 0.895 3.835 0.895 3.835 0.775 3.955 0.775 3.955 0.815 3.965 0.815 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.575 0.72 3.54 0.72 3.54 1.04 3.46 1.04 3.46 0.725 3.395 0.725 3.395 0.64 3.575 0.64 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.405 0.895 0.315 0.895 0.315 1.025 0.235 1.025 0.235 0.895 0.23 0.895 0.23 0.775 0.325 0.775 0.325 0.62 0.405 0.62 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.125 0.335 1.125 0.335 1.65 1.385 1.65 1.385 1.54 1.505 1.54 1.505 1.65 2.295 1.65 2.295 1.25 2.415 1.25 2.415 1.31 2.355 1.31 2.355 1.65 3.175 1.65 3.175 1.41 3.295 1.41 3.295 1.47 3.235 1.47 3.235 1.65 4.03 1.65 4.03 0.995 4.09 0.995 4.09 1.65 4.46 1.65 4.46 1.025 4.52 1.025 4.52 1.65 4.885 1.65 4.885 0.965 4.945 0.965 4.945 1.65 5.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 0.06 5.05 0.06 5.05 0.17 4.93 0.17 4.93 0.06 4.55 0.06 4.55 0.2 4.49 0.2 4.49 0.06 4.09 0.06 4.09 0.17 3.97 0.17 3.97 0.06 3.415 0.06 3.415 0.17 3.295 0.17 3.295 0.06 2.415 0.06 2.415 0.47 2.355 0.47 2.355 0.06 1.505 0.06 1.505 0.17 1.385 0.17 1.385 0.06 0.305 0.06 0.305 0.275 0.365 0.275 0.365 0.335 0.245 0.335 0.245 0.06 0 0.06 0 -0.06 5.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.285 0.565 5.18 0.565 5.18 1.085 5.12 1.085 5.12 0.725 4.84 0.725 4.84 0.665 5.12 0.665 5.12 0.505 5.285 0.505 ;
      POLYGON 5.27 0.38 4.525 0.38 4.525 0.925 4.395 0.925 4.395 0.805 4.465 0.805 4.465 0.38 4.125 0.38 4.125 0.635 4.135 0.635 4.135 0.755 4.065 0.755 4.065 0.38 2.635 0.38 2.635 0.93 2.695 0.93 2.695 0.99 2.575 0.99 2.575 0.63 2.315 0.63 2.315 0.68 2.195 0.68 2.195 0.62 2.255 0.62 2.255 0.57 2.575 0.57 2.575 0.32 5.27 0.32 ;
      POLYGON 3.855 0.54 3.735 0.54 3.735 1.09 3.76 1.09 3.76 1.15 3.64 1.15 3.64 1.09 3.675 1.09 3.675 0.54 3.295 0.54 3.295 0.83 3.175 0.83 3.175 0.48 3.855 0.48 ;
      POLYGON 3.035 0.54 2.855 0.54 2.855 1.03 2.9 1.03 2.9 1.15 0.865 1.15 0.865 0.97 0.725 0.97 0.725 0.52 0.665 0.52 0.665 0.46 0.785 0.46 0.785 0.91 0.925 0.91 0.925 1.09 2.795 1.09 2.795 0.48 3.035 0.48 ;
      POLYGON 2.475 0.99 1.855 0.99 1.855 0.43 1.915 0.43 1.915 0.93 2.415 0.93 2.415 0.73 2.475 0.73 ;
      POLYGON 2.135 0.83 2.015 0.83 2.015 0.33 0.945 0.33 0.945 0.75 1.02 0.75 1.02 0.81 0.885 0.81 0.885 0.33 0.565 0.33 0.565 1.09 0.54 1.09 0.54 1.15 0.48 1.15 0.48 1.03 0.505 1.03 0.505 0.39 0.485 0.39 0.485 0.27 1.785 0.27 1.785 0.17 1.905 0.17 1.905 0.27 2.075 0.27 2.075 0.77 2.135 0.77 ;
      RECT 1.12 1.25 1.94 1.33 ;
      POLYGON 1.755 0.99 1.635 0.99 1.635 0.63 1.37 0.63 1.37 0.72 1.31 0.72 1.31 0.57 1.62 0.57 1.62 0.46 1.74 0.46 1.74 0.52 1.695 0.52 1.695 0.93 1.755 0.93 ;
      POLYGON 1.535 0.88 1.18 0.88 1.18 0.99 1.04 0.99 1.04 0.93 1.12 0.93 1.12 0.52 1.045 0.52 1.045 0.46 1.18 0.46 1.18 0.82 1.475 0.82 1.475 0.73 1.535 0.73 ;
      POLYGON 0.405 0.52 0.13 0.52 0.13 1.15 0.07 1.15 0.07 0.27 0.13 0.27 0.13 0.46 0.405 0.46 ;
  END
END EDFFX2

MACRO EDFFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFX4 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6938 LAYER Metal1 ;
    ANTENNADIFFAREA 4.02455 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4554 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.111111 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 63.5177865 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.715 1.44 5.655 1.44 5.655 1.11 5.305 1.11 5.305 1.44 5.245 1.44 5.245 1.05 5.26 1.05 5.26 0.63 5.1 0.63 5.1 0.57 5.69 0.57 5.69 0.63 5.32 0.63 5.32 0.98 5.34 0.98 5.34 1.05 5.715 1.05 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6938 LAYER Metal1 ;
    ANTENNADIFFAREA 4.02455 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4554 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.111111 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 63.5177865 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.895 1.44 4.835 1.44 4.835 1.11 4.485 1.11 4.485 1.44 4.425 1.44 4.425 1.05 4.46 1.05 4.46 0.63 4.16 0.63 4.16 0.57 4.75 0.57 4.75 0.63 4.52 0.63 4.52 0.98 4.54 0.98 4.54 1.05 4.895 1.05 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.645 0.815 4.145 0.895 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.165 1.115 3.045 1.115 3.045 0.895 2.885 0.895 2.885 0.815 3.165 0.815 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.765 0.34 1.265 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 1.77 0 1.77 0 1.65 0.395 1.65 0.395 1.36 0.455 1.36 0.455 1.65 1.5 1.65 1.5 1.185 1.62 1.185 1.62 1.245 1.56 1.245 1.56 1.65 2.49 1.65 2.49 1.49 2.61 1.49 2.61 1.55 2.55 1.55 2.55 1.65 2.96 1.65 2.96 1.49 3.08 1.49 3.08 1.55 3.02 1.55 3.02 1.65 4.2 1.65 4.2 1.32 4.26 1.32 4.26 1.65 4.63 1.65 4.63 1.21 4.69 1.21 4.69 1.65 5.04 1.65 5.04 1.05 5.1 1.05 5.1 1.65 5.45 1.65 5.45 1.21 5.51 1.21 5.51 1.65 5.88 1.65 5.88 1.08 5.94 1.08 5.94 1.65 6.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 0.06 6.01 0.06 6.01 0.52 5.95 0.52 5.95 0.06 5.455 0.06 5.455 0.17 5.335 0.17 5.335 0.06 4.985 0.06 4.985 0.17 4.865 0.17 4.865 0.06 4.515 0.06 4.515 0.17 4.395 0.17 4.395 0.06 4.045 0.06 4.045 0.17 3.925 0.17 3.925 0.06 2.99 0.06 2.99 0.555 2.93 0.555 2.93 0.06 2.55 0.06 2.55 0.465 2.61 0.465 2.61 0.525 2.49 0.525 2.49 0.06 1.56 0.06 1.56 0.19 1.62 0.19 1.62 0.25 1.5 0.25 1.5 0.06 0.425 0.06 0.425 0.505 0.365 0.505 0.365 0.06 0 0.06 0 -0.06 6.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.215 1.44 6.085 1.44 6.085 0.98 5.815 0.98 5.815 0.78 5.875 0.78 5.875 0.92 6.155 0.92 6.155 0.54 6.215 0.54 ;
      POLYGON 6.055 0.82 5.995 0.82 5.995 0.68 5.79 0.68 5.79 0.47 4.91 0.47 4.91 0.85 4.77 0.85 4.77 0.79 4.85 0.79 4.85 0.47 3.58 0.47 3.58 0.555 3.52 0.555 3.52 0.39 3.15 0.39 3.15 0.715 2.785 0.715 2.785 1.09 2.845 1.09 2.845 1.15 2.725 1.15 2.725 0.77 2.405 0.77 2.405 0.71 2.725 0.71 2.725 0.52 2.785 0.52 2.785 0.655 3.09 0.655 3.09 0.33 3.58 0.33 3.58 0.41 5.85 0.41 5.85 0.62 6.055 0.62 ;
      POLYGON 4.325 1.075 3.73 1.075 3.73 1.18 3.65 1.18 3.65 0.995 4.245 0.995 4.245 0.815 4.325 0.815 ;
      POLYGON 4.055 1.235 3.89 1.235 3.89 1.34 3.55 1.34 3.55 1.435 3.275 1.435 3.275 1.375 3.49 1.375 3.49 1.055 3.485 1.055 3.485 0.715 3.425 0.715 3.425 0.655 3.68 0.655 3.68 0.57 3.88 0.57 3.88 0.63 3.74 0.63 3.74 0.715 3.545 0.715 3.545 0.995 3.55 0.995 3.55 1.28 3.83 1.28 3.83 1.175 4.055 1.175 ;
      POLYGON 3.405 0.55 3.325 0.55 3.325 1.155 3.39 1.155 3.39 1.275 3.175 1.275 3.175 1.34 1.72 1.34 1.72 1.085 1.4 1.085 1.4 1.34 0.975 1.34 0.975 1.215 0.8 1.215 0.8 0.505 0.86 0.505 0.86 1.155 1.035 1.155 1.035 1.28 1.34 1.28 1.34 1.025 1.78 1.025 1.78 1.28 3.115 1.28 3.115 1.215 3.265 1.215 3.265 0.49 3.405 0.49 ;
      POLYGON 2.625 1.12 2.195 1.12 2.195 1.15 2.075 1.15 2.075 1.09 2.085 1.09 2.085 0.505 2.145 0.505 2.145 1.06 2.565 1.06 2.565 0.87 2.625 0.87 ;
      POLYGON 2.305 0.96 2.245 0.96 2.245 0.405 1.78 0.405 1.78 0.41 1.34 0.41 1.34 0.405 1.02 0.405 1.02 0.87 1.08 0.87 1.08 0.93 0.96 0.93 0.96 0.405 0.66 0.405 0.66 1.385 0.6 1.385 0.6 0.345 1.23 0.345 1.23 0.295 1.35 0.295 1.35 0.345 1.4 0.345 1.4 0.35 1.72 0.35 1.72 0.345 1.98 0.345 1.98 0.295 2.1 0.295 2.1 0.345 2.305 0.345 ;
      POLYGON 1.94 1.18 1.88 1.18 1.88 0.765 1.395 0.765 1.395 0.705 1.88 0.705 1.88 0.505 1.94 0.505 ;
      POLYGON 1.725 0.925 1.24 0.925 1.24 1.18 1.18 1.18 1.18 0.595 1.12 0.595 1.12 0.535 1.24 0.535 1.24 0.865 1.725 0.865 ;
      POLYGON 0.5 0.745 0.44 0.745 0.44 0.665 0.16 0.665 0.16 1.36 0.205 1.36 0.205 1.48 0.145 1.48 0.145 1.42 0.1 1.42 0.1 0.605 0.16 0.605 0.16 0.41 0.22 0.41 0.22 0.605 0.5 0.605 ;
  END
END EDFFX4

MACRO EDFFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN EDFFXL 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.969825 LAYER Metal1 ;
    ANTENNADIFFAREA 3.1169 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2106 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.10173325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 108.66096875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.54 1.145 5.46 1.145 5.46 0.79 5.47 0.79 5.47 0.415 5.54 0.415 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.930125 LAYER Metal1 ;
    ANTENNADIFFAREA 3.1169 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2106 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.913224 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 107.83475775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.54 0.8 4.53 0.8 4.53 1.02 4.45 1.02 4.45 0.75 4.46 0.75 4.46 0.65 4.42 0.65 4.42 0.57 4.54 0.57 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 20.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.14 0.92 4.1 0.92 4.1 1.32 3.495 1.32 3.495 1.465 3.17 1.465 3.17 1.405 3.435 1.405 3.435 0.705 3.495 0.705 3.495 1.26 4.04 1.26 4.04 0.86 4.06 0.86 4.06 0.79 4.14 0.79 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.765 0.755 3.94 1.16 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.765 0.34 1.265 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 0 1.77 0 1.65 0.395 1.65 0.395 1.36 0.455 1.36 0.455 1.65 1.675 1.65 1.675 1.52 1.615 1.52 1.615 1.46 1.735 1.46 1.735 1.65 2.815 1.65 2.815 1.51 2.875 1.51 2.875 1.65 3.87 1.65 3.87 1.42 3.99 1.42 3.99 1.48 3.93 1.48 3.93 1.65 4.685 1.65 4.685 0.995 4.745 0.995 4.745 1.65 5.215 1.65 5.215 1.12 5.275 1.12 5.275 1.65 5.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5.26 0.06 5.26 0.51 5.2 0.51 5.2 0.06 4.775 0.06 4.775 0.2 4.715 0.2 4.715 0.06 3.93 0.06 3.93 0.215 3.99 0.215 3.99 0.275 3.87 0.275 3.87 0.06 2.815 0.06 2.815 0.54 2.875 0.54 2.875 0.6 2.755 0.6 2.755 0.06 1.675 0.06 1.675 0.225 1.735 0.225 1.735 0.285 1.615 0.285 1.615 0.06 0.425 0.06 0.425 0.505 0.365 0.505 0.365 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.37 0.69 5 0.69 5 1.02 4.92 1.02 4.92 0.66 4.88 0.66 4.88 0.54 4.96 0.54 4.96 0.58 5 0.58 5 0.61 5.37 0.61 ;
      POLYGON 4.615 0.435 3.13 0.435 3.13 1.085 3.16 1.085 3.16 1.145 3.04 1.145 3.04 0.985 2.74 0.985 2.74 0.865 2.8 0.865 2.8 0.925 3.07 0.925 3.07 0.375 4.615 0.375 ;
      POLYGON 4.32 1.13 4.2 1.13 4.2 1.07 4.26 1.07 4.26 0.655 3.665 0.655 3.665 0.99 3.605 0.99 3.605 0.595 4.25 0.595 4.25 0.535 4.31 0.535 4.31 0.595 4.32 0.595 ;
      POLYGON 3.335 1.305 2.675 1.305 2.675 1.36 2.295 1.36 2.295 1.28 1.995 1.28 1.995 1.2 1.355 1.2 1.355 1.28 0.815 1.28 0.815 0.535 0.875 0.535 0.875 1.22 1.295 1.22 1.295 1.14 2.055 1.14 2.055 1.22 2.355 1.22 2.355 1.3 2.615 1.3 2.615 1.245 3.275 1.245 3.275 0.535 3.335 0.535 ;
      POLYGON 2.97 0.825 2.91 0.825 2.91 0.76 2.64 0.76 2.64 1.14 2.515 1.14 2.515 1.2 2.455 1.2 2.455 1.08 2.58 1.08 2.58 0.76 2.475 0.76 2.475 0.535 2.535 0.535 2.535 0.7 2.97 0.7 ;
      POLYGON 2.48 0.98 2.42 0.98 2.42 0.92 2.315 0.92 2.315 0.825 2.155 0.825 2.155 0.705 2.315 0.705 2.315 0.445 1.455 0.445 1.455 0.435 1.035 0.435 1.035 0.955 0.975 0.955 0.975 0.435 0.66 0.435 0.66 1.385 0.6 1.385 0.6 0.375 1.2 0.375 1.2 0.275 1.32 0.275 1.32 0.375 1.515 0.375 1.515 0.385 2.375 0.385 2.375 0.86 2.48 0.86 ;
      POLYGON 2.275 1.12 2.155 1.12 2.155 0.985 1.52 0.985 1.52 0.9 1.995 0.9 1.995 0.545 2.115 0.545 2.115 0.605 2.055 0.605 2.055 0.925 2.215 0.925 2.215 1.06 2.275 1.06 ;
      POLYGON 2.195 1.44 1.835 1.44 1.835 1.36 1.515 1.36 1.515 1.44 1.15 1.44 1.15 1.38 1.455 1.38 1.455 1.3 1.895 1.3 1.895 1.38 2.195 1.38 ;
      POLYGON 1.84 0.795 1.195 0.795 1.195 1.12 1.02 1.12 1.02 1.06 1.135 1.06 1.135 0.565 1.255 0.565 1.255 0.625 1.195 0.625 1.195 0.735 1.84 0.735 ;
      POLYGON 0.5 0.775 0.44 0.775 0.44 0.665 0.16 0.665 0.16 1.36 0.205 1.36 0.205 1.48 0.145 1.48 0.145 1.42 0.1 1.42 0.1 0.605 0.16 0.605 0.16 0.41 0.22 0.41 0.22 0.605 0.5 0.605 ;
  END
END EDFFXL

MACRO FILL1
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILL1 0 0 ;
  SIZE 0.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 0.2 1.77 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 0.2 0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END FILL1

MACRO FILL16
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILL16 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 3.2 1.77 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 3.2 0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END FILL16

MACRO FILL2
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILL2 0 0 ;
  SIZE 0.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 0.4 1.77 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 0.4 0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END FILL2

MACRO FILL32
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILL32 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 6.4 1.77 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 6.4 0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END FILL32

MACRO FILL4
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILL4 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 0.8 1.77 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 0.8 0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END FILL4

MACRO FILL64
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILL64 0 0 ;
  SIZE 12.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 12.8 1.77 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 12.8 0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END FILL64

MACRO FILL8
  CLASS CORE SPACER ;
  ORIGIN 0 0 ;
  FOREIGN FILL8 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 1.6 1.77 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 1.6 0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END FILL8

MACRO FSWNX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FSWNX1 0 0 ;
  SIZE 6.2 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN ExtVSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "ExtVSS ExtVSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.235 2.34 4.965 2.34 4.965 3.12 0.68 3.12 0.68 2.01 0.74 2.01 0.74 2.92 1.09 2.92 1.09 2.01 1.15 2.01 1.15 2.92 1.5 2.92 1.5 2.01 1.56 2.01 1.56 2.92 1.91 2.92 1.91 2.01 1.97 2.01 1.97 2.92 2.32 2.92 2.32 2.01 2.38 2.01 2.38 2.92 2.73 2.92 2.73 2.01 2.79 2.01 2.79 2.92 3.14 2.92 3.14 2.01 3.2 2.01 3.2 2.92 3.55 2.92 3.55 2.01 3.61 2.01 3.61 2.92 3.96 2.92 3.96 2.01 4.02 2.01 4.02 2.92 4.37 2.92 4.37 2.01 4.43 2.01 4.43 2.92 4.765 2.92 4.765 2.28 5.175 2.28 5.175 2.05 5.235 2.05 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.645 1.54 4.765 1.54 4.765 0.5 4.43 0.5 4.43 1.41 4.37 1.41 4.37 0.5 4.02 0.5 4.02 1.41 3.96 1.41 3.96 0.5 3.61 0.5 3.61 1.41 3.55 1.41 3.55 0.5 3.2 0.5 3.2 1.41 3.14 1.41 3.14 0.5 2.79 0.5 2.79 1.41 2.73 1.41 2.73 0.5 2.38 0.5 2.38 1.41 2.32 1.41 2.32 0.5 1.97 0.5 1.97 1.41 1.91 1.41 1.91 0.5 1.56 0.5 1.56 1.41 1.5 1.41 1.5 0.5 1.15 0.5 1.15 1.41 1.09 1.41 1.09 0.5 0.74 0.5 0.74 1.41 0.68 1.41 0.68 0.3 4.965 0.3 4.965 0.775 4.825 0.775 4.825 1.48 5.175 1.48 5.175 1.11 5.235 1.11 5.235 1.48 5.585 1.48 5.585 1.11 5.645 1.11 ;
    END
  END ExtVSS
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 4.635 1.77 4.635 2.81 4.575 2.81 4.575 1.86 4.225 1.86 4.225 2.81 4.165 2.81 4.165 1.86 3.815 1.86 3.815 2.81 3.755 2.81 3.755 1.86 3.405 1.86 3.405 2.81 3.345 2.81 3.345 1.86 2.995 1.86 2.995 2.81 2.935 2.81 2.935 1.86 2.585 1.86 2.585 2.81 2.525 2.81 2.525 1.86 2.175 1.86 2.175 2.81 2.115 2.81 2.115 1.86 1.765 1.86 1.765 2.81 1.705 2.81 1.705 1.86 1.355 1.86 1.355 2.81 1.295 2.81 1.295 1.86 0.945 1.86 0.945 2.81 0.885 2.81 0.885 1.86 0.535 1.86 0.535 2.81 0.475 2.81 0.475 1.77 0 1.77 0 1.65 0.475 1.65 0.475 0.61 0.535 0.61 0.535 1.56 0.885 1.56 0.885 0.61 0.945 0.61 0.945 1.56 1.295 1.56 1.295 0.61 1.355 0.61 1.355 1.56 1.705 1.56 1.705 0.61 1.765 0.61 1.765 1.56 2.115 1.56 2.115 0.61 2.175 0.61 2.175 1.56 2.525 1.56 2.525 0.61 2.585 0.61 2.585 1.56 2.935 1.56 2.935 0.61 2.995 0.61 2.995 1.56 3.345 1.56 3.345 0.61 3.405 0.61 3.405 1.56 3.755 1.56 3.755 0.61 3.815 0.61 3.815 1.56 4.165 1.56 4.165 0.61 4.225 0.61 4.225 1.56 4.575 1.56 4.575 0.61 4.635 0.61 4.635 1.65 6.2 1.65 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 3.48 0 3.48 0 3.36 5.175 3.36 5.175 2.7 5.235 2.7 5.235 3.36 6.2 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 5.645 0.06 5.645 0.72 5.585 0.72 5.585 0.06 5.235 0.06 5.235 0.72 5.175 0.72 5.175 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
  END VDD
  PIN PSOn_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.83995 LAYER Metal1 ;
    ANTENNADIFFAREA 7.0771 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.17675 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.66237525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 39.7323135 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.85 2.585 5.44 2.585 5.44 3.09 5.38 3.09 5.38 2.05 5.44 2.05 5.44 2.43 5.85 2.43 ;
    END
  END PSOn_out
  PIN PSOn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.98 0.83 6.145 0.99 ;
    END
  END PSOn
  OBS
    LAYER Metal1 ;
      POLYGON 5.88 1.395 5.82 1.395 5.82 0.94 5.525 0.94 5.525 0.88 5.82 0.88 5.82 0.32 5.88 0.32 ;
      POLYGON 5.44 1.41 5.38 1.41 5.38 0.94 5.005 0.94 5.005 1.36 4.945 1.36 4.945 0.88 5.38 0.88 5.38 0.27 5.44 0.27 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END FSWNX1

MACRO FSWX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FSWX1 0 0 ;
  SIZE 6.2 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN ExtVSS
    DIRECTION INOUT ;
    USE GROUND ;
    NETEXPR "ExtVSS ExtVSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.645 1.54 4.765 1.54 4.765 0.5 4.43 0.5 4.43 1.41 4.37 1.41 4.37 0.5 4.02 0.5 4.02 1.41 3.96 1.41 3.96 0.5 3.61 0.5 3.61 1.41 3.55 1.41 3.55 0.5 3.2 0.5 3.2 1.41 3.14 1.41 3.14 0.5 2.79 0.5 2.79 1.41 2.73 1.41 2.73 0.5 2.38 0.5 2.38 1.41 2.32 1.41 2.32 0.5 1.97 0.5 1.97 1.41 1.91 1.41 1.91 0.5 1.56 0.5 1.56 1.41 1.5 1.41 1.5 0.5 1.15 0.5 1.15 1.41 1.09 1.41 1.09 0.5 0.74 0.5 0.74 1.41 0.68 1.41 0.68 0.3 4.965 0.3 4.965 0.715 4.825 0.715 4.825 1.48 5.175 1.48 5.175 1.11 5.235 1.11 5.235 1.48 5.585 1.48 5.585 1.11 5.645 1.11 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6.055 2.31 5.995 2.31 5.995 1.94 5.645 1.94 5.645 2.31 5.585 2.31 5.585 1.94 5.235 1.94 5.235 2.31 5.175 2.31 5.175 1.94 4.965 1.94 4.965 3.12 0.68 3.12 0.68 2.01 0.74 2.01 0.74 2.92 1.09 2.92 1.09 2.01 1.15 2.01 1.15 2.92 1.5 2.92 1.5 2.01 1.56 2.01 1.56 2.92 1.91 2.92 1.91 2.01 1.97 2.01 1.97 2.92 2.32 2.92 2.32 2.01 2.38 2.01 2.38 2.92 2.73 2.92 2.73 2.01 2.79 2.01 2.79 2.92 3.14 2.92 3.14 2.01 3.2 2.01 3.2 2.92 3.55 2.92 3.55 2.01 3.61 2.01 3.61 2.92 3.96 2.92 3.96 2.01 4.02 2.01 4.02 2.92 4.37 2.92 4.37 2.01 4.43 2.01 4.43 2.92 4.765 2.92 4.765 1.88 6.055 1.88 ;
    END
  END ExtVSS
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 4.635 1.77 4.635 2.81 4.575 2.81 4.575 1.86 4.225 1.86 4.225 2.81 4.165 2.81 4.165 1.86 3.815 1.86 3.815 2.81 3.755 2.81 3.755 1.86 3.405 1.86 3.405 2.81 3.345 2.81 3.345 1.86 2.995 1.86 2.995 2.81 2.935 2.81 2.935 1.86 2.585 1.86 2.585 2.81 2.525 2.81 2.525 1.86 2.175 1.86 2.175 2.81 2.115 2.81 2.115 1.86 1.765 1.86 1.765 2.81 1.705 2.81 1.705 1.86 1.355 1.86 1.355 2.81 1.295 2.81 1.295 1.86 0.945 1.86 0.945 2.81 0.885 2.81 0.885 1.86 0.535 1.86 0.535 2.81 0.475 2.81 0.475 1.77 0 1.77 0 1.65 0.475 1.65 0.475 0.61 0.535 0.61 0.535 1.56 0.885 1.56 0.885 0.61 0.945 0.61 0.945 1.56 1.295 1.56 1.295 0.61 1.355 0.61 1.355 1.56 1.705 1.56 1.705 0.61 1.765 0.61 1.765 1.56 2.115 1.56 2.115 0.61 2.175 0.61 2.175 1.56 2.525 1.56 2.525 0.61 2.585 0.61 2.585 1.56 2.935 1.56 2.935 0.61 2.995 0.61 2.995 1.56 3.345 1.56 3.345 0.61 3.405 0.61 3.405 1.56 3.755 1.56 3.755 0.61 3.815 0.61 3.815 1.56 4.165 1.56 4.165 0.61 4.225 0.61 4.225 1.56 4.575 1.56 4.575 0.61 4.635 0.61 4.635 1.65 6.2 1.65 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 3.48 0 3.48 0 3.36 5.175 3.36 5.175 2.7 5.235 2.7 5.235 3.36 5.585 3.36 5.585 2.7 5.645 2.7 5.645 3.36 5.995 3.36 5.995 2.7 6.055 2.7 6.055 3.36 6.2 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 5.645 0.06 5.645 0.72 5.585 0.72 5.585 0.06 5.235 0.06 5.235 0.72 5.175 0.72 5.175 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
  END VDD
  PIN PSO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.088889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.535 0.85 5.885 0.97 ;
    END
  END PSO
  PIN PSO_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.0528 LAYER Metal1 ;
    ANTENNADIFFAREA 7.5576 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.215 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.627819 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 39.99753075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.85 3.15 5.79 3.15 5.79 2.56 5.44 2.56 5.44 3.15 5.38 3.15 5.38 2.01 5.44 2.01 5.44 2.46 5.79 2.46 5.79 2.01 5.85 2.01 ;
    END
  END PSO_out
  OBS
    LAYER Metal1 ;
      POLYGON 5.44 1.41 5.38 1.41 5.38 0.94 5.065 0.94 5.065 1.36 5.005 1.36 5.005 0.88 5.38 0.88 5.38 0.27 5.44 0.27 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END FSWX1

MACRO HOLDX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HOLDX1 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3495 LAYER Metal1 ;
    ANTENNADIFFAREA 0.57745 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.07785 LAYER Metal1 ;
      ANTENNAMAXAREACAR 4.48940275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 36.49325625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 1.02 0.87 1.02 0.87 0.98 0.34 0.98 0.34 0.74 0.4 0.74 0.4 0.92 0.86 0.92 0.86 0.79 0.87 0.79 0.87 0.54 0.94 0.54 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.435 1.65 0.435 1.275 0.495 1.275 0.495 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.495 0.06 0.495 0.2 0.435 0.2 0.435 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.58 0.82 0.52 0.82 0.52 0.64 0.24 0.64 0.24 1.29 0.18 1.29 0.18 0.52 0.26 0.52 0.26 0.58 0.58 0.58 ;
  END
END HOLDX1

MACRO HSWDNX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HSWDNX1 0 0 ;
  SIZE 6.2 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.3 3.2 2.635 3.2 2.635 2.65 1.845 2.65 1.845 1.97 1.665 1.97 1.665 2.495 1.605 2.495 1.605 1.97 1.255 1.97 1.255 2.495 1.195 2.495 1.195 1.97 0.81 1.97 0.81 2.495 0.75 2.495 0.75 1.97 0.66 1.97 0.66 1.91 1.905 1.91 1.905 2.59 2.44 2.59 2.44 1.89 2.5 1.89 2.5 2.59 2.635 2.59 2.635 1.87 2.885 1.87 2.885 3.015 3.19 3.015 3.19 1.9 3.25 1.9 3.25 3.015 3.6 3.015 3.6 1.9 3.66 1.9 3.66 3.015 4.01 3.015 4.01 1.9 4.07 1.9 4.07 3.015 4.42 3.015 4.42 1.9 4.48 1.9 4.48 3.015 4.83 3.015 4.83 1.9 4.89 1.9 4.89 3.015 5.24 3.015 5.24 1.9 5.3 1.9 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.3 1.52 5.24 1.52 5.24 0.375 4.89 0.375 4.89 1.52 4.83 1.52 4.83 0.375 4.48 0.375 4.48 1.52 4.42 1.52 4.42 0.375 4.07 0.375 4.07 1.52 4.01 1.52 4.01 0.375 3.66 0.375 3.66 1.52 3.6 1.52 3.6 0.375 3.25 0.375 3.25 1.52 3.19 1.52 3.19 0.375 2.88 0.375 2.88 1.52 0.66 1.52 0.66 1.46 0.75 1.46 0.75 0.9 0.81 0.9 0.81 1.46 1.16 1.46 1.16 0.9 1.22 0.9 1.22 1.46 1.57 1.46 1.57 0.9 1.63 0.9 1.63 1.46 1.89 1.46 1.89 0.905 1.95 0.905 1.95 1.46 2.3 1.46 2.3 0.905 2.36 0.905 2.36 1.46 2.63 1.46 2.63 0.19 5.3 0.19 ;
    END
  END ExtVDD
  PIN PSO1n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.135 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.0444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.605 0.625 0.89 0.81 ;
    END
  END PSO1n
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 3.48 0 3.48 0 3.36 0.75 3.36 0.75 2.795 0.81 2.795 0.81 3.36 1.195 3.36 1.195 2.795 1.255 2.795 1.255 3.36 1.605 3.36 1.605 2.795 1.665 2.795 1.665 3.36 6.2 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 2.28 0.06 2.28 0.6 2.22 0.6 2.22 0.06 1.87 0.06 1.87 0.6 1.81 0.6 1.81 0.06 1.63 0.06 1.63 0.545 1.57 0.545 1.57 0.06 1.22 0.06 1.22 0.545 1.16 0.545 1.16 0.06 0.81 0.06 0.81 0.545 0.75 0.545 0.75 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 5.095 1.77 5.095 2.92 5.035 2.92 5.035 1.77 4.685 1.77 4.685 2.92 4.625 2.92 4.625 1.77 4.275 1.77 4.275 2.92 4.215 2.92 4.215 1.77 3.865 1.77 3.865 2.92 3.805 2.92 3.805 1.77 3.455 1.77 3.455 2.92 3.395 2.92 3.395 1.77 3.045 1.77 3.045 2.92 2.985 2.92 2.985 1.77 2.11 1.77 2.11 2.495 2.05 2.495 2.05 1.77 0 1.77 0 1.65 2.985 1.65 2.985 0.5 3.045 0.5 3.045 1.65 3.395 1.65 3.395 0.5 3.455 0.5 3.455 1.65 3.805 1.65 3.805 0.5 3.865 0.5 3.865 1.65 4.215 1.65 4.215 0.5 4.275 0.5 4.275 1.65 4.625 1.65 4.625 0.5 4.685 0.5 4.685 1.65 5.035 1.65 5.035 0.5 5.095 0.5 5.095 1.65 6.2 1.65 ;
    END
  END VDD
  PIN PSO2n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.03375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.73333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.88 2.675 0.41 2.675 0.41 2.5 0.62 2.5 0.62 2.555 0.88 2.555 ;
    END
  END PSO2n
  PIN PSO1n_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.751025 LAYER Metal1 ;
    ANTENNADIFFAREA 6.9195 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.12725 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.98893325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 40.63339975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.195 0.92 2.155 0.92 2.155 1.355 2.095 1.355 2.095 0.92 2.065 0.92 2.065 0.79 2.095 0.79 2.095 0.66 2.015 0.66 2.015 0.3 2.075 0.3 2.075 0.6 2.155 0.6 2.155 0.79 2.195 0.79 ;
    END
  END PSO1n_out
  PIN PSO2n_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.676975 LAYER Metal1 ;
    ANTENNADIFFAREA 6.87 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.12725 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.9232425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 40.31536925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.53 2.44 1.46 2.44 1.46 3.095 1.4 3.095 1.4 2.44 1.385 2.44 1.385 2.31 1.4 2.31 1.4 2.045 1.46 2.045 1.46 2.31 1.53 2.31 ;
    END
  END PSO2n_out
  OBS
    LAYER Metal1 ;
      POLYGON 1.79 1.295 1.73 1.295 1.73 0.76 1.425 0.76 1.425 1.35 1.365 1.35 1.365 0.76 1.015 0.76 1.015 1.35 0.955 1.35 0.955 0.245 1.015 0.245 1.015 0.7 1.365 0.7 1.365 0.245 1.425 0.245 1.425 0.7 1.73 0.7 1.73 0.695 1.79 0.695 ;
      POLYGON 1.3 2.675 1.015 2.675 1.015 3.095 0.955 3.095 0.955 2.045 1.015 2.045 1.015 2.615 1.3 2.615 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END HSWDNX1

MACRO HSWDX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HSWDX1 0 0 ;
  SIZE 6.4 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN PSO1_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.63595 LAYER Metal1 ;
    ANTENNADIFFAREA 7.0436 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.2195 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.4415335 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 38.7466175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.665 0.225 2.725 1.35 ;
    END
  END PSO1_out
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.62 3.2 2.95 3.2 2.95 2.6 2.185 2.6 2.185 1.93 1.8 1.93 1.8 2.465 1.74 2.465 1.74 1.93 1.345 1.93 1.345 2.465 1.285 2.465 1.285 1.93 0.9 1.93 0.9 2.405 0.84 2.405 0.84 1.87 1.095 1.87 1.095 1.85 1.215 1.85 1.215 1.87 2.245 1.87 2.245 2.54 2.66 2.54 2.66 1.995 2.72 1.995 2.72 2.54 2.95 2.54 2.95 1.87 3.07 1.87 3.07 3.015 3.42 3.015 3.42 1.9 3.48 1.9 3.48 3.015 3.83 3.015 3.83 1.9 3.89 1.9 3.89 3.015 4.24 3.015 4.24 1.9 4.3 1.9 4.3 3.015 4.65 3.015 4.65 1.9 4.71 1.9 4.71 3.015 5.06 3.015 5.06 1.9 5.12 1.9 5.12 3.015 5.47 3.015 5.47 1.9 5.53 1.9 5.53 3.015 5.62 3.015 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.63 0.375 5.53 0.375 5.53 1.52 5.47 1.52 5.47 0.375 5.12 0.375 5.12 1.52 5.06 1.52 5.06 0.375 4.71 0.375 4.71 1.52 4.65 1.52 4.65 0.375 4.3 0.375 4.3 1.52 4.24 1.52 4.24 0.375 3.89 0.375 3.89 1.52 3.83 1.52 3.83 0.375 3.48 0.375 3.48 1.52 3.42 1.52 3.42 0.375 3.07 0.375 3.07 1.52 0.835 1.52 0.835 0.9 0.895 0.9 0.895 1.46 1.28 1.46 1.28 0.9 1.34 0.9 1.34 1.46 1.69 1.46 1.69 0.9 1.75 0.9 1.75 1.46 2.1 1.46 2.1 0.9 2.16 0.9 2.16 1.46 2.46 1.46 2.46 0.96 2.52 0.96 2.52 1.46 2.95 1.46 2.95 0.19 5.63 0.19 ;
    END
  END ExtVDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 3.48 0 3.48 0 3.36 0.835 3.36 0.835 3.02 0.84 3.02 0.84 2.82 0.9 2.82 0.9 3.08 0.895 3.08 0.895 3.36 1.285 3.36 1.285 2.82 1.345 2.82 1.345 3.36 1.74 3.36 1.74 2.82 1.8 2.82 1.8 3.36 6.4 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 0.06 2.52 0.06 2.52 0.485 2.46 0.485 2.46 0.06 2.16 0.06 2.16 0.525 2.1 0.525 2.1 0.06 1.75 0.06 1.75 0.525 1.69 0.525 1.69 0.06 1.34 0.06 1.34 0.525 1.28 0.525 1.28 0.06 0.895 0.06 0.895 0.485 0.835 0.485 0.835 0.06 0 0.06 0 -0.06 6.4 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 1.77 5.325 1.77 5.325 2.92 5.265 2.92 5.265 1.77 4.915 1.77 4.915 2.92 4.855 2.92 4.855 1.77 4.505 1.77 4.505 2.92 4.445 2.92 4.445 1.77 4.095 1.77 4.095 2.92 4.035 2.92 4.035 1.77 3.685 1.77 3.685 2.92 3.625 2.92 3.625 1.77 3.275 1.77 3.275 2.92 3.215 2.92 3.215 1.77 2.45 1.77 2.45 2.465 2.39 2.465 2.39 1.77 0 1.77 0 1.65 3.215 1.65 3.215 0.5 3.275 0.5 3.275 1.65 3.625 1.65 3.625 0.5 3.685 0.5 3.685 1.65 4.035 1.65 4.035 0.5 4.095 0.5 4.095 1.65 4.445 1.65 4.445 0.5 4.505 0.5 4.505 1.65 4.855 1.65 4.855 0.5 4.915 0.5 4.915 1.65 5.265 1.65 5.265 0.5 5.325 0.5 5.325 1.65 6.4 1.65 ;
    END
  END VDD
  PIN PSO2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.17948725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.965 2.7 0.66 2.7 0.66 2.5 0.795 2.5 0.795 2.58 0.965 2.58 ;
    END
  END PSO2
  PIN PSO1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.4358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.97 0.695 0.965 0.695 0.965 0.785 0.835 0.785 0.835 0.585 0.965 0.585 0.965 0.635 0.97 0.635 ;
    END
  END PSO1
  PIN PSO2_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.70345 LAYER Metal1 ;
    ANTENNADIFFAREA 6.9716 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.2195 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.496884 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 39.0381305 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.165 3.01 2.005 3.01 2.005 3.08 1.945 3.08 1.945 2.075 2.005 2.075 2.005 2.715 2.165 2.715 ;
    END
  END PSO2_out
  OBS
    LAYER Metal1 ;
      POLYGON 2.33 1.135 2.27 1.135 2.27 1.115 2.26 1.115 2.26 0.775 1.955 0.775 1.955 1.35 1.895 1.35 1.895 0.775 1.545 0.775 1.545 1.35 1.485 1.35 1.485 0.225 1.545 0.225 1.545 0.715 1.895 0.715 1.895 0.225 1.955 0.225 1.955 0.715 2.32 0.715 2.32 0.895 2.33 0.895 ;
      POLYGON 1.59 3.3 1.49 3.3 1.49 2.015 1.55 2.015 1.55 3.18 1.59 3.18 ;
      POLYGON 1.415 0.755 1.235 0.755 1.235 0.695 1.1 0.695 1.1 1.29 1.04 1.29 1.04 0.225 1.1 0.225 1.1 0.635 1.415 0.635 ;
      POLYGON 1.395 2.665 1.105 2.665 1.105 3.08 1.045 3.08 1.045 2.015 1.105 2.015 1.105 2.605 1.395 2.605 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END HSWDX1

MACRO HSWNX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HSWNX1 0 0 ;
  SIZE 7.2 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.385 3.25 2.105 3.25 2.105 1.93 2.005 1.93 2.005 2.41 1.945 2.41 1.945 1.93 1.325 1.93 1.325 2.485 1.265 2.485 1.265 1.93 0.915 1.93 0.915 2.485 0.855 2.485 0.855 1.93 0.68 1.93 0.68 1.87 2.165 1.87 2.165 1.845 2.225 1.845 2.225 3.025 2.575 3.025 2.575 1.845 2.635 1.845 2.635 3.025 2.985 3.025 2.985 1.845 3.045 1.845 3.045 3.025 3.395 3.025 3.395 1.845 3.455 1.845 3.455 3.025 3.805 3.025 3.805 1.845 3.865 1.845 3.865 3.025 4.215 3.025 4.215 1.845 4.275 1.845 4.275 3.025 4.625 3.025 4.625 1.845 4.685 1.845 4.685 3.025 5.035 3.025 5.035 1.845 5.095 1.845 5.095 3.025 5.445 3.025 5.445 1.845 5.505 1.845 5.505 3.025 5.855 3.025 5.855 1.845 5.915 1.845 5.915 3.025 6.265 3.025 6.265 1.845 6.385 1.845 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6.385 1.545 6.325 1.545 6.325 1.575 6.265 1.575 6.265 0.395 5.915 0.395 5.915 1.575 5.855 1.575 5.855 0.395 5.505 0.395 5.505 1.575 5.445 1.575 5.445 0.395 5.095 0.395 5.095 1.575 5.035 1.575 5.035 0.395 4.685 0.395 4.685 1.575 4.625 1.575 4.625 0.395 4.275 0.395 4.275 1.575 4.215 1.575 4.215 0.395 3.865 0.395 3.865 1.575 3.805 1.575 3.805 0.395 3.455 0.395 3.455 1.575 3.395 1.575 3.395 0.395 3.045 0.395 3.045 1.575 2.985 1.575 2.985 0.395 2.635 0.395 2.635 1.575 2.575 1.575 2.575 0.395 2.225 0.395 2.225 1.575 2.165 1.575 2.165 1.55 0.68 1.55 0.68 1.49 0.755 1.49 0.755 1.42 0.75 1.42 0.75 0.97 0.81 0.97 0.81 1.35 0.815 1.35 0.815 1.49 1.16 1.49 1.16 0.97 1.22 0.97 1.22 1.49 1.57 1.49 1.57 0.97 1.63 0.97 1.63 1.49 1.94 1.49 1.94 1.015 2 1.015 2 1.49 2.105 1.49 2.105 0.17 6.385 0.17 ;
    END
  END ExtVDD
  PIN PSOn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.911111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.97 2.715 0.78 2.715 0.78 2.82 0.635 2.82 0.635 2.5 0.78 2.5 0.78 2.595 0.97 2.595 ;
    END
  END PSOn
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 3.48 0 3.48 0 3.36 0.855 3.36 0.855 2.82 0.915 2.82 0.915 3.36 1.265 3.36 1.265 2.82 1.325 2.82 1.325 3.36 7.2 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 0.06 1.63 0.06 1.63 0.555 1.57 0.555 1.57 0.06 1.22 0.06 1.22 0.555 1.16 0.555 1.16 0.06 0.815 0.06 0.815 0.36 0.81 0.36 0.81 0.555 0.75 0.555 0.75 0.255 0.755 0.255 0.755 0.06 0 0.06 0 -0.06 7.2 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 1.77 6.12 1.77 6.12 2.865 6.06 2.865 6.06 1.77 5.71 1.77 5.71 2.865 5.65 2.865 5.65 1.77 5.3 1.77 5.3 2.865 5.24 2.865 5.24 1.77 4.89 1.77 4.89 2.865 4.83 2.865 4.83 1.77 4.48 1.77 4.48 2.865 4.42 2.865 4.42 1.77 4.07 1.77 4.07 2.865 4.01 2.865 4.01 1.77 3.66 1.77 3.66 2.865 3.6 2.865 3.6 1.77 3.25 1.77 3.25 2.865 3.19 2.865 3.19 1.77 2.84 1.77 2.84 2.865 2.78 2.865 2.78 1.77 2.43 1.77 2.43 2.865 2.37 2.865 2.37 1.77 0 1.77 0 1.65 2.37 1.65 2.37 0.555 2.43 0.555 2.43 1.65 2.78 1.65 2.78 0.555 2.84 0.555 2.84 1.65 3.19 1.65 3.19 0.555 3.25 0.555 3.25 1.65 3.6 1.65 3.6 0.555 3.66 0.555 3.66 1.65 4.01 1.65 4.01 0.555 4.07 0.555 4.07 1.65 4.42 1.65 4.42 0.555 4.48 0.555 4.48 1.65 4.83 1.65 4.83 0.555 4.89 0.555 4.89 1.65 5.24 1.65 5.24 0.555 5.3 0.555 5.3 1.65 5.65 1.65 5.65 0.555 5.71 0.555 5.71 1.65 6.06 1.65 6.06 0.555 6.12 0.555 6.12 1.65 7.2 1.65 ;
    END
  END VDD
  PIN PSOn_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.529675 LAYER Metal1 ;
    ANTENNADIFFAREA 8.8632 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.7955 LAYER Metal1 ;
      ANTENNAMAXAREACAR 4.75058475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 31.06599825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.425 1.42 1.365 1.42 1.365 0.735 1.015 0.735 1.015 1.42 0.955 1.42 0.955 0.255 1.015 0.255 1.015 0.625 1.365 0.625 1.365 0.255 1.425 0.255 ;
    END
  END PSOn_out
  OBS
    LAYER Metal1 ;
      POLYGON 1.81 2.685 1.12 2.685 1.12 3.12 1.06 3.12 1.06 2.035 1.12 2.035 1.12 2.625 1.75 2.625 1.75 2.065 1.81 2.065 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END HSWNX1

MACRO HSWX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HSWX1 0 0 ;
  SIZE 7.2 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.365 3.25 1.805 3.25 1.805 3.025 1.925 3.025 1.925 1.945 1.64 1.945 1.64 1.98 1.59 1.98 1.59 2.48 1.53 2.48 1.53 1.98 1.46 1.98 1.46 1.945 1.37 1.945 1.37 2.48 1.31 2.48 1.31 1.945 0.96 1.945 0.96 2.48 0.9 2.48 0.9 1.885 1.46 1.885 1.46 1.86 1.64 1.86 1.64 1.885 1.985 1.885 1.985 1.845 2.045 1.845 2.045 3.025 2.395 3.025 2.395 1.845 2.455 1.845 2.455 3.025 2.805 3.025 2.805 1.845 2.865 1.845 2.865 3.025 3.215 3.025 3.215 1.845 3.275 1.845 3.275 3.025 3.625 3.025 3.625 1.845 3.685 1.845 3.685 3.025 4.035 3.025 4.035 1.845 4.095 1.845 4.095 3.025 4.445 3.025 4.445 1.845 4.505 1.845 4.505 3.025 4.855 3.025 4.855 1.845 4.915 1.845 4.915 3.025 5.265 3.025 5.265 1.845 5.325 1.845 5.325 3.025 5.675 3.025 5.675 1.845 5.735 1.845 5.735 3.025 6.085 3.025 6.085 1.845 6.145 1.845 6.145 3.025 6.305 3.025 6.305 1.905 6.365 1.905 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6.365 1.53 6.305 1.53 6.305 0.395 6.145 0.395 6.145 1.58 6.085 1.58 6.085 0.395 5.735 0.395 5.735 1.575 5.675 1.575 5.675 0.395 5.325 0.395 5.325 1.575 5.265 1.575 5.265 0.395 4.915 0.395 4.915 1.575 4.855 1.575 4.855 0.395 4.505 0.395 4.505 1.575 4.445 1.575 4.445 0.395 4.095 0.395 4.095 1.575 4.035 1.575 4.035 0.395 3.685 0.395 3.685 1.575 3.625 1.575 3.625 0.395 3.275 0.395 3.275 1.575 3.215 1.575 3.215 0.395 2.865 0.395 2.865 1.575 2.805 1.575 2.805 0.395 2.455 0.395 2.455 1.575 2.395 1.575 2.395 0.395 2.045 0.395 2.045 1.575 1.985 1.575 1.985 1.545 1.64 1.545 1.64 1.575 1.46 1.575 1.46 1.545 1.11 1.545 1.11 0.935 1.17 0.935 1.17 1.485 1.46 1.485 1.46 1.455 1.535 1.455 1.535 0.935 1.595 0.935 1.595 1.455 1.64 1.455 1.64 1.485 1.925 1.485 1.925 0.395 1.815 0.395 1.815 0.17 6.365 0.17 ;
    END
  END ExtVDD
  PIN PSO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.28205125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 0.6 1.165 0.79 ;
    END
  END PSO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 3.48 0 3.48 0 3.36 0.9 3.36 0.9 2.82 0.96 2.82 0.96 3.36 1.31 3.36 1.31 2.82 1.37 2.82 1.37 3.36 7.2 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 0.06 1.17 0.06 1.17 0.535 1.11 0.535 1.11 0.06 0 0.06 0 -0.06 7.2 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 1.77 5.94 1.77 5.94 2.865 5.88 2.865 5.88 1.77 5.53 1.77 5.53 2.865 5.47 2.865 5.47 1.77 5.12 1.77 5.12 2.865 5.06 2.865 5.06 1.77 4.71 1.77 4.71 2.865 4.65 2.865 4.65 1.77 4.3 1.77 4.3 2.865 4.24 2.865 4.24 1.77 3.89 1.77 3.89 2.865 3.83 2.865 3.83 1.77 3.48 1.77 3.48 2.865 3.42 2.865 3.42 1.77 3.07 1.77 3.07 2.865 3.01 2.865 3.01 1.77 2.66 1.77 2.66 2.865 2.6 2.865 2.6 1.77 2.25 1.77 2.25 2.865 2.19 2.865 2.19 1.77 0 1.77 0 1.65 2.19 1.65 2.19 0.555 2.25 0.555 2.25 1.65 2.6 1.65 2.6 0.555 2.66 0.555 2.66 1.65 3.01 1.65 3.01 0.555 3.07 0.555 3.07 1.65 3.42 1.65 3.42 0.555 3.48 0.555 3.48 1.65 3.83 1.65 3.83 0.555 3.89 0.555 3.89 1.65 4.24 1.65 4.24 0.555 4.3 0.555 4.3 1.65 4.65 1.65 4.65 0.555 4.71 0.555 4.71 1.65 5.06 1.65 5.06 0.555 5.12 0.555 5.12 1.65 5.47 1.65 5.47 0.555 5.53 0.555 5.53 1.65 5.88 1.65 5.88 0.555 5.94 0.555 5.94 1.65 7.2 1.65 ;
    END
  END VDD
  PIN PSO_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.445 LAYER Metal1 ;
    ANTENNADIFFAREA 8.7862 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.75725 LAYER Metal1 ;
      ANTENNAMAXAREACAR 4.8058045 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 31.52539475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.57 0.54 1.375 0.54 1.375 1.325 1.315 1.325 1.315 0.275 1.375 0.275 1.375 0.41 1.57 0.41 ;
    END
  END PSO_out
  OBS
    LAYER Metal1 ;
      POLYGON 1.855 2.72 1.165 2.72 1.165 3.12 1.105 3.12 1.105 2.03 1.165 2.03 1.165 2.66 1.855 2.66 ;
      POLYGON 0.965 1.545 0.845 1.545 0.845 1.485 0.905 1.485 0.905 0.275 0.965 0.275 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END HSWX1

MACRO INVX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX1 0 0 ;
  SIZE 0.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1734 LAYER Metal1 ;
    ANTENNADIFFAREA 0.34455 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.33 1.29 0.27 1.29 0.27 0.8 0.25 0.8 0.25 0.68 0.27 0.68 0.27 0.37 0.33 0.37 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.05 0.59 0.19 0.8 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.4 1.77 0 1.77 0 1.65 0.08 1.65 0.08 1.46 0.14 1.46 0.14 1.65 0.4 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.4 0.06 0.14 0.06 0.14 0.2 0.08 0.2 0.08 0.06 0 0.06 0 -0.06 0.4 -0.06 ;
    END
  END VSS
END INVX1

MACRO INVX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX12 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9636 LAYER Metal1 ;
    ANTENNADIFFAREA 1.9176 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.18 0.8 2.1 0.8 2.1 0.77 1.975 0.77 1.975 1.37 1.915 1.37 1.915 0.96 1.565 0.96 1.565 1.37 1.505 1.37 1.505 0.96 1.155 0.96 1.155 1.37 1.095 1.37 1.095 0.96 0.745 0.96 0.745 1.37 0.685 1.37 0.685 0.96 0.335 0.96 0.335 1.37 0.275 1.37 0.275 0.96 0.27 0.96 0.27 0.9 1.915 0.9 1.915 0.69 0.275 0.69 0.275 0.35 0.335 0.35 0.335 0.63 0.685 0.63 0.685 0.35 0.745 0.35 0.745 0.63 1.095 0.63 1.095 0.35 1.155 0.35 1.155 0.63 1.505 0.63 1.505 0.35 1.565 0.35 1.565 0.63 1.915 0.63 1.915 0.35 1.975 0.35 1.975 0.705 2.18 0.705 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.351 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.6068375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.82 0.215 0.82 0.215 0.87 0.07 0.87 0.07 0.72 0.215 0.72 0.215 0.76 1.8 0.76 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 0.06 2.18 0.06 2.18 0.63 2.12 0.63 2.12 0.06 1.77 0.06 1.77 0.47 1.71 0.47 1.71 0.06 1.36 0.06 1.36 0.47 1.3 0.47 1.3 0.06 0.95 0.06 0.95 0.47 0.89 0.47 0.89 0.06 0.54 0.06 0.54 0.47 0.48 0.47 0.48 0.06 0.13 0.06 0.13 0.66 0.07 0.66 0.07 0.06 0 0.06 0 -0.06 2.4 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.935 0.13 0.935 0.13 1.65 0.48 1.65 0.48 1.095 0.54 1.095 0.54 1.65 0.89 1.65 0.89 1.095 0.95 1.095 0.95 1.65 1.3 1.65 1.3 1.095 1.36 1.095 1.36 1.65 1.71 1.65 1.71 1.095 1.77 1.095 1.77 1.65 2.12 1.65 2.12 0.935 2.18 0.935 2.18 1.65 2.4 1.65 ;
    END
  END VDD
END INVX12

MACRO INVX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX16 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2858 LAYER Metal1 ;
    ANTENNADIFFAREA 2.5144 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 0.8 2.92 0.8 2.92 0.77 2.795 0.77 2.795 1.345 2.735 1.345 2.735 0.96 2.385 0.96 2.385 1.345 2.325 1.345 2.325 0.96 1.975 0.96 1.975 1.345 1.915 1.345 1.915 0.96 1.565 0.96 1.565 1.345 1.505 1.345 1.505 0.96 1.155 0.96 1.155 1.345 1.095 1.345 1.095 0.96 0.745 0.96 0.745 1.345 0.685 1.345 0.685 0.96 0.335 0.96 0.335 1.345 0.275 1.345 0.275 0.9 2.735 0.9 2.735 0.69 0.275 0.69 0.275 0.365 0.335 0.365 0.335 0.63 0.685 0.63 0.685 0.365 0.745 0.365 0.745 0.63 1.095 0.63 1.095 0.365 1.155 0.365 1.155 0.63 1.505 0.63 1.505 0.365 1.565 0.365 1.565 0.63 1.915 0.63 1.915 0.365 1.975 0.365 1.975 0.63 2.325 0.63 2.325 0.365 2.385 0.365 2.385 0.63 2.735 0.63 2.735 0.365 2.795 0.365 2.795 0.705 3 0.705 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4662 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.73745175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.62 0.82 0.215 0.82 0.215 0.87 0.07 0.87 0.07 0.72 0.215 0.72 0.215 0.76 2.62 0.76 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 0.06 3 0.06 3 0.63 2.94 0.63 2.94 0.06 2.59 0.06 2.59 0.485 2.53 0.485 2.53 0.06 2.18 0.06 2.18 0.485 2.12 0.485 2.12 0.06 1.77 0.06 1.77 0.485 1.71 0.485 1.71 0.06 1.36 0.06 1.36 0.485 1.3 0.485 1.3 0.06 0.95 0.06 0.95 0.485 0.89 0.485 0.89 0.06 0.54 0.06 0.54 0.485 0.48 0.485 0.48 0.06 0.13 0.06 0.13 0.66 0.07 0.66 0.07 0.06 0 0.06 0 -0.06 3.2 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.935 0.13 0.935 0.13 1.65 0.48 1.65 0.48 1.07 0.54 1.07 0.54 1.65 0.89 1.65 0.89 1.07 0.95 1.07 0.95 1.65 1.3 1.65 1.3 1.07 1.36 1.07 1.36 1.65 1.71 1.65 1.71 1.07 1.77 1.07 1.77 1.65 2.12 1.65 2.12 1.07 2.18 1.07 2.18 1.65 2.53 1.65 2.53 1.07 2.59 1.07 2.59 1.65 2.94 1.65 2.94 0.935 3 0.935 3 1.65 3.2 1.65 ;
    END
  END VDD
END INVX16

MACRO INVX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX2 0 0 ;
  SIZE 0.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2663 LAYER Metal1 ;
    ANTENNADIFFAREA 0.48725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.53 0.8 0.335 0.8 0.335 1.29 0.265 1.29 0.265 0.4 0.335 0.4 0.335 0.72 0.53 0.72 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.79487175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.045 0.6 0.195 0.8 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 0.06 0.53 0.06 0.53 0.64 0.47 0.64 0.47 0.06 0.17 0.06 0.17 0.21 0.045 0.21 0.045 0.06 0 0.06 0 -0.06 0.6 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 1.77 0 1.77 0 1.65 0.045 1.65 0.045 1.46 0.17 1.46 0.17 1.65 0.47 1.65 0.47 0.9 0.53 0.9 0.53 1.65 0.6 1.65 ;
    END
  END VDD
END INVX2

MACRO INVX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX20 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2419 LAYER Metal1 ;
    ANTENNADIFFAREA 3.0846 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.615 1.36 3.555 1.36 3.555 0.96 3.205 0.96 3.205 1.36 3.145 1.36 3.145 0.96 2.795 0.96 2.795 1.36 2.735 1.36 2.735 0.96 2.385 0.96 2.385 1.36 2.325 1.36 2.325 0.96 1.975 0.96 1.975 1.36 1.915 1.36 1.915 0.96 1.565 0.96 1.565 1.36 1.505 1.36 1.505 0.96 1.155 0.96 1.155 1.36 1.095 1.36 1.095 0.96 0.745 0.96 0.745 1.36 0.685 1.36 0.685 0.96 0.335 0.96 0.335 1.36 0.275 1.36 0.275 0.9 3.535 0.9 3.535 0.69 0.275 0.69 0.275 0.355 0.335 0.355 0.335 0.63 0.685 0.63 0.685 0.355 0.745 0.355 0.745 0.63 1.095 0.63 1.095 0.355 1.155 0.355 1.155 0.63 1.505 0.63 1.505 0.355 1.565 0.355 1.565 0.63 1.915 0.63 1.915 0.355 1.975 0.355 1.975 0.63 2.325 0.63 2.325 0.355 2.385 0.355 2.385 0.63 2.735 0.63 2.735 0.355 2.795 0.355 2.795 0.63 3.145 0.63 3.145 0.355 3.205 0.355 3.205 0.63 3.555 0.63 3.555 0.355 3.615 0.355 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.585225 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.801871 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.435 0.82 0.215 0.82 0.215 0.87 0.07 0.87 0.07 0.72 0.215 0.72 0.215 0.76 3.435 0.76 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 0.06 3.41 0.06 3.41 0.475 3.35 0.475 3.35 0.06 3 0.06 3 0.475 2.94 0.475 2.94 0.06 2.59 0.06 2.59 0.475 2.53 0.475 2.53 0.06 2.18 0.06 2.18 0.475 2.12 0.475 2.12 0.06 1.77 0.06 1.77 0.475 1.71 0.475 1.71 0.06 1.36 0.06 1.36 0.475 1.3 0.475 1.3 0.06 0.95 0.06 0.95 0.475 0.89 0.475 0.89 0.06 0.54 0.06 0.54 0.475 0.48 0.475 0.48 0.06 0.13 0.06 0.13 0.66 0.07 0.66 0.07 0.06 0 0.06 0 -0.06 3.8 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.935 0.13 0.935 0.13 1.65 0.48 1.65 0.48 1.085 0.54 1.085 0.54 1.65 0.89 1.65 0.89 1.085 0.95 1.085 0.95 1.65 1.3 1.65 1.3 1.085 1.36 1.085 1.36 1.65 1.71 1.65 1.71 1.085 1.77 1.085 1.77 1.65 2.12 1.65 2.12 1.085 2.18 1.085 2.18 1.65 2.53 1.65 2.53 1.085 2.59 1.085 2.59 1.65 2.94 1.65 2.94 1.085 3 1.085 3 1.65 3.35 1.65 3.35 1.11 3.41 1.11 3.41 1.65 3.8 1.65 ;
    END
  END VDD
END INVX20

MACRO INVX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX3 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3169 LAYER Metal1 ;
    ANTENNADIFFAREA 0.64145 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.73 1.29 0.67 1.29 0.67 0.8 0.32 0.8 0.32 1.29 0.26 1.29 0.26 0.4 0.32 0.4 0.32 0.72 0.67 0.72 0.67 0.4 0.73 0.4 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.08775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.12820525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.055 0.62 0.16 0.845 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 0.06 0.525 0.06 0.525 0.66 0.465 0.66 0.465 0.06 0.17 0.06 0.17 0.21 0.04 0.21 0.04 0.06 0 0.06 0 -0.06 0.8 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.77 0 1.77 0 1.65 0.04 1.65 0.04 1.46 0.17 1.46 0.17 1.65 0.465 1.65 0.465 0.905 0.525 0.905 0.525 1.65 0.8 1.65 ;
    END
  END VDD
END INVX3

MACRO INVX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX4 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4191 LAYER Metal1 ;
    ANTENNADIFFAREA 0.78365 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.95 0.935 0.745 0.935 0.745 1.34 0.685 1.34 0.685 0.94 0.335 0.94 0.335 1.34 0.275 1.34 0.275 0.875 0.87 0.875 0.87 0.695 0.275 0.695 0.275 0.395 0.335 0.395 0.335 0.63 0.685 0.63 0.685 0.395 0.745 0.395 0.745 0.625 0.95 0.625 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.20512825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.785 0.815 0.215 0.815 0.215 0.865 0.07 0.865 0.07 0.72 0.215 0.72 0.215 0.755 0.785 0.755 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.96 0.06 0.96 0.22 0.825 0.22 0.825 0.06 0.54 0.06 0.54 0.515 0.48 0.515 0.48 0.06 0.13 0.06 0.13 0.655 0.07 0.655 0.07 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.95 0.13 0.95 0.13 1.65 0.48 1.65 0.48 1.09 0.54 1.09 0.54 1.65 0.825 1.65 0.825 1.51 0.96 1.51 0.96 1.65 1 1.65 ;
    END
  END VDD
END INVX4

MACRO INVX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX6 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5319 LAYER Metal1 ;
    ANTENNADIFFAREA 1.0536 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.155 1.37 1.095 1.37 1.095 0.94 0.745 0.94 0.745 1.37 0.685 1.37 0.685 0.94 0.335 0.94 0.335 1.37 0.275 1.37 0.275 0.88 1.075 0.88 1.075 0.69 0.275 0.69 0.275 0.35 0.335 0.35 0.335 0.63 0.685 0.63 0.685 0.35 0.745 0.35 0.745 0.63 1.095 0.63 1.095 0.35 1.155 0.35 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.72649575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.98 0.82 0.07 0.82 0.07 0.72 0.15 0.72 0.15 0.76 0.98 0.76 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.935 0.13 0.935 0.13 1.65 0.48 1.65 0.48 1.085 0.54 1.085 0.54 1.65 0.89 1.65 0.89 1.085 0.95 1.085 0.95 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 0.95 0.06 0.95 0.47 0.89 0.47 0.89 0.06 0.54 0.06 0.54 0.47 0.48 0.47 0.48 0.06 0.13 0.06 0.13 0.66 0.07 0.66 0.07 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END INVX6

MACRO INVX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX8 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.02845 LAYER Metal1 ;
    ANTENNADIFFAREA 1.3496 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.565 1.345 1.505 1.345 1.505 0.94 1.155 0.94 1.155 1.345 1.095 1.345 1.095 0.94 0.745 0.94 0.745 1.345 0.685 1.345 0.685 0.94 0.335 0.94 0.335 1.345 0.275 1.345 0.275 0.88 1.485 0.88 1.485 0.7 0.275 0.7 0.275 0.365 0.335 0.365 0.335 0.635 0.685 0.635 0.685 0.365 0.745 0.365 0.745 0.63 1.095 0.63 1.095 0.365 1.155 0.365 1.155 0.63 1.505 0.63 1.505 0.365 1.565 0.365 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.82110675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.385 0.82 0.07 0.82 0.07 0.72 0.15 0.72 0.15 0.76 1.385 0.76 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.935 0.13 0.935 0.13 1.65 0.48 1.65 0.48 1.095 0.54 1.095 0.54 1.65 0.89 1.65 0.89 1.095 0.95 1.095 0.95 1.65 1.3 1.65 1.3 1.095 1.36 1.095 1.36 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.36 0.06 1.36 0.485 1.3 0.485 1.3 0.06 0.95 0.06 0.95 0.485 0.89 0.485 0.89 0.06 0.54 0.06 0.54 0.485 0.48 0.485 0.48 0.06 0.13 0.06 0.13 0.66 0.07 0.66 0.07 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END INVX8

MACRO INVXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVXL 0 0 ;
  SIZE 0.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.190875 LAYER Metal1 ;
    ANTENNADIFFAREA 0.241025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.27 0.405 0.35 1.205 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.055 0.59 0.17 0.8 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.4 0.06 0.145 0.06 0.145 0.21 0.085 0.21 0.085 0.06 0 0.06 0 -0.06 0.4 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.4 1.77 0 1.77 0 1.65 0.055 1.65 0.055 1.475 0.18 1.475 0.18 1.65 0.4 1.65 ;
    END
  END VDD
END INVXL

MACRO ISOHLDX1_OFF
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ISOHLDX1_OFF 0 0 ;
  SIZE 3.6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 3.6 1.77 ;
    END
  END VDD
  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 0.74 1.19 0.92 ;
    END
  END ISO
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0176 LAYER Metal1 ;
    ANTENNADIFFAREA 1.654 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1395 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.4630825 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 115.2903225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.965 2.63 2.775 2.63 2.775 3.16 2.715 3.16 2.715 2.07 2.775 2.07 2.775 2.5 2.965 2.5 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.63 0.6 2.765 0.8 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 3.48 0 3.48 0 3.36 1.49 3.36 1.49 2.965 1.55 2.965 1.55 3.36 2.51 3.36 2.51 2.9 2.57 2.9 2.57 3.36 3.6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 0.06 2.76 0.06 2.76 0.455 2.7 0.455 2.7 0.06 1.655 0.06 1.655 0.46 1.595 0.46 1.595 0.06 0 0.06 0 -0.06 3.6 -0.06 ;
    END
  END VSS
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.57 2.46 2.51 2.46 2.51 1.93 1.55 1.93 1.55 2.325 1.49 2.325 1.49 1.93 0.95 1.93 0.95 2.49 1.055 2.49 1.055 2.61 0.755 2.61 0.755 2.49 0.89 2.49 0.89 1.87 2.57 1.87 ;
    END
  END ExtVDD
  OBS
    LAYER Metal1 ;
      POLYGON 2.76 1.525 1.135 1.525 1.135 1.465 1.595 1.465 1.595 1.075 1.655 1.075 1.655 1.465 2.7 1.465 2.7 1.09 2.76 1.09 ;
      POLYGON 2.65 2.77 2.365 2.77 2.365 3.16 2.305 3.16 2.305 2.07 2.365 2.07 2.365 2.71 2.65 2.71 ;
      POLYGON 2.45 1.305 2.39 1.305 2.39 1.23 1.985 1.23 1.985 1.17 2.39 1.17 2.39 0.31 2.45 0.31 ;
      POLYGON 2.24 0.94 2.22 0.94 2.22 0.965 2.16 0.965 2.16 0.94 1.86 0.94 1.86 1.29 1.8 1.29 1.8 0.88 2.16 0.88 2.16 0.46 1.78 0.46 1.78 0.4 1.8 0.4 1.8 0.315 1.86 0.315 1.86 0.4 2.22 0.4 2.22 0.88 2.24 0.88 ;
      POLYGON 2.14 2.865 1.86 2.865 1.86 3.11 1.8 3.11 1.8 2.865 1.445 2.865 1.445 2.895 1.385 2.895 1.385 2.415 1.445 2.415 1.445 2.805 2.08 2.805 2.08 2.325 1.8 2.325 1.8 2.11 1.86 2.11 1.86 2.265 2.14 2.265 ;
      POLYGON 1.99 2.715 1.565 2.715 1.565 2.595 1.625 2.595 1.625 2.655 1.99 2.655 ;
      POLYGON 1.75 0.675 1.45 0.675 1.45 1.29 1.39 1.29 1.39 0.315 1.45 0.315 1.45 0.615 1.75 0.615 ;
      POLYGON 1.345 2.325 1.26 2.325 1.26 2.625 1.32 2.625 1.32 2.685 1.26 2.685 1.26 2.965 1.345 2.965 1.345 3.11 1.285 3.11 1.285 3.025 1.2 3.025 1.2 2.265 1.285 2.265 1.285 2.11 1.345 2.11 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END ISOHLDX1_OFF

MACRO ISOHLDX1_ON
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ISOHLDX1_ON 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.77 0 1.77 0 1.65 0.355 1.65 0.355 1.275 0.415 1.275 0.415 1.65 1.11 1.65 1.11 1.275 1.41 1.275 1.41 1.65 2.125 1.65 2.125 1.275 2.185 1.275 2.185 1.65 2.57 1.65 2.57 1.1 2.63 1.1 2.63 1.65 3 1.65 ;
    END
  END VDD
  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.83333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.98 0.445 1.11 ;
    END
  END ISO
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.74845 LAYER Metal1 ;
    ANTENNADIFFAREA 1.5303 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1395 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.53369175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 90.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.97 1.11 2.835 1.11 2.835 1.49 2.775 1.49 2.775 0.21 2.835 0.21 2.835 0.98 2.97 0.98 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 17.4074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.165 0.515 1.14 0.515 1.14 0.73 1.095 0.73 1.095 1.215 1.035 1.215 1.035 0.485 1.015 0.485 1.015 0.425 1.165 0.425 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 0.06 2.63 0.06 2.63 0.47 2.57 0.47 2.57 0.06 2.185 0.06 2.185 0.355 2.125 0.355 2.125 0.06 1.41 0.06 1.41 0.355 1.11 0.355 1.11 0.06 0.415 0.06 0.415 0.355 0.355 0.355 0.355 0.06 0 0.06 0 -0.06 3 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.705 0.925 2.425 0.925 2.425 1.49 2.365 1.49 2.365 0.21 2.425 0.21 2.425 0.865 2.705 0.865 ;
      POLYGON 1.935 1.19 1.875 1.19 1.875 1.49 1.815 1.49 1.815 1.13 1.875 1.13 1.875 0.505 1.815 0.505 1.815 0.21 1.875 0.21 1.875 0.445 1.935 0.445 ;
      POLYGON 1.78 0.925 1.615 0.925 1.615 1.49 1.555 1.49 1.555 0.21 1.615 0.21 1.615 0.865 1.78 0.865 ;
      RECT 1.69 0.395 1.75 0.785 ;
      RECT 1.275 0.415 1.335 1.205 ;
      RECT 0.8 0.21 0.86 1.49 ;
      POLYGON 0.71 0.755 0.62 0.755 0.62 1.06 0.71 1.06 0.71 1.12 0.62 1.12 0.62 1.49 0.56 1.49 0.56 0.21 0.62 0.21 0.62 0.695 0.71 0.695 ;
      POLYGON 0.495 0.795 0.465 0.795 0.465 0.8 0.405 0.8 0.405 0.795 0.2 0.795 0.2 1.275 0.21 1.275 0.21 1.49 0.15 1.49 0.15 1.355 0.14 1.355 0.14 0.735 0.15 0.735 0.15 0.21 0.21 0.21 0.21 0.735 0.495 0.735 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END ISOHLDX1_ON

MACRO ISOHX1_OFF
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ISOHX1_OFF 0 0 ;
  SIZE 2.8 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6945 LAYER Metal1 ;
    ANTENNADIFFAREA 0.6981 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 23.74358975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 193.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.885 1.95 1.945 3.18 ;
    END
  END Y
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 2.58 1.605 2.58 1.605 2.61 1.305 2.61 1.305 1.93 0.83 1.93 0.83 2.265 0.77 2.265 0.77 1.87 1.365 1.87 1.365 2.49 1.605 2.49 1.605 2.52 1.68 2.52 1.68 1.95 1.74 1.95 ;
    END
  END ExtVDD
  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.83333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.815 2.675 1.01 2.795 ;
    END
  END ISO
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.388889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.56 2.425 0.785 2.545 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 3.48 0 3.48 0 3.36 0.63 3.36 0.63 3.005 0.69 3.005 0.69 3.36 1.04 3.36 1.04 3.005 1.1 3.005 1.1 3.36 1.68 3.36 1.68 2.92 1.74 2.92 1.74 3.36 2.8 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 2.8 0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT -0.005 1.65 2.8 1.77 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.825 2.79 1.14 2.79 1.14 2.935 0.895 2.935 0.895 3.15 0.835 3.15 0.835 2.875 1.08 2.875 1.08 2.05 1.14 2.05 1.14 2.73 1.825 2.73 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END ISOHX1_OFF

MACRO ISOHX1_ON
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ISOHX1_ON 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.175 1.65 0.175 1.14 0.235 1.14 0.235 1.65 0.725 1.65 0.725 1.025 0.785 1.025 0.785 1.65 1.2 1.65 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.16 0.59 0.34 0.74 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4953 LAYER Metal1 ;
    ANTENNADIFFAREA 0.59385 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.93333325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 139.64102575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.99 1.415 0.93 1.415 0.93 1.11 0.86 1.11 0.86 0.98 0.93 0.98 0.93 0.24 0.99 0.24 ;
    END
  END Y
  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.5555555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.41 0.77 0.54 0.94 ;
    END
  END ISO
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.785 0.06 0.785 0.5 0.725 0.5 0.725 0.06 0.345 0.06 0.345 0.445 0.285 0.445 0.285 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.87 0.855 0.665 0.855 0.665 1.17 0.545 1.17 0.545 1.355 0.485 1.355 0.485 1.11 0.605 1.11 0.605 0.565 0.49 0.565 0.49 0.3 0.55 0.3 0.55 0.505 0.665 0.505 0.665 0.795 0.87 0.795 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END ISOHX1_ON

MACRO ISOLX1_OFF
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ISOLX1_OFF 0 0 ;
  SIZE 2.8 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2453 LAYER Metal1 ;
    ANTENNADIFFAREA 1.1419 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXAREACAR 27.39934 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 204.02640275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.89 1.95 1.95 3.18 ;
    END
  END Y
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.745 2.58 1.61 2.58 1.61 2.61 1.31 2.61 1.31 2.575 1.16 2.575 1.16 1.94 0.81 1.94 0.81 2.265 0.75 2.265 0.75 1.88 1.22 1.88 1.22 2.515 1.31 2.515 1.31 2.49 1.61 2.49 1.61 2.52 1.685 2.52 1.685 2.01 1.485 2.01 1.485 1.95 1.745 1.95 ;
    END
  END ExtVDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.555 2.485 0.86 2.605 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 3.48 0 3.48 0 3.36 1.045 3.36 1.045 3.005 1.105 3.005 1.105 3.36 1.685 3.36 1.685 2.92 1.745 2.92 1.745 3.36 2.8 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 0.06 1.275 0.06 1.275 0.47 1.215 0.47 1.215 0.06 0 0.06 0 -0.06 2.8 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 2.8 1.77 ;
    END
  END VDD
  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.12962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.145 0.625 1.41 0.745 ;
    END
  END ISO
  OBS
    LAYER Metal1 ;
      POLYGON 1.83 2.79 1.015 2.79 1.015 2.795 0.795 2.795 0.795 3.15 0.735 3.15 0.735 2.735 0.955 2.735 0.955 2.05 1.015 2.05 1.015 2.73 1.83 2.73 ;
      POLYGON 1.605 1.345 1.215 1.345 1.215 0.93 1.275 0.93 1.275 1.285 1.605 1.285 ;
      RECT 1.01 0.325 1.07 1.54 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END ISOLX1_OFF

MACRO ISOLX1_ON
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ISOLX1_ON 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6798 LAYER Metal1 ;
    ANTENNADIFFAREA 0.7303 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.95709575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 126.5346535 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 0.92 1.275 0.92 1.275 1.475 1.215 1.475 1.215 0.235 1.275 0.235 1.275 0.79 1.365 0.79 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.115 1.65 0.115 1.26 0.175 1.26 0.175 1.65 0.57 1.65 0.57 1.26 0.63 1.26 0.63 1.65 1.01 1.65 1.01 1.085 1.07 1.085 1.07 1.65 1.4 1.65 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.92 0.675 1.11 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 1.07 0.06 1.07 0.495 1.01 0.495 1.01 0.06 0.175 0.06 0.175 0.38 0.115 0.38 0.115 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
  END VSS
  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.31481475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.03 0.595 0.22 0.8 ;
    END
  END ISO
  OBS
    LAYER Metal1 ;
      POLYGON 1.145 0.985 0.835 0.985 0.835 1.475 0.775 1.475 0.775 0.925 1.025 0.925 1.025 0.64 0.67 0.64 0.67 0.29 0.73 0.29 0.73 0.58 1.085 0.58 1.085 0.925 1.145 0.925 ;
      POLYGON 0.92 0.805 0.38 0.805 0.38 1.475 0.32 1.475 0.32 0.235 0.38 0.235 0.38 0.745 0.92 0.745 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END ISOLX1_ON

MACRO ISONLX1_OFF
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ISONLX1_OFF 0 0 ;
  SIZE 2.8 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6903 LAYER Metal1 ;
    ANTENNADIFFAREA 0.7051 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 23.6 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 191.79487175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.89 1.95 1.95 3.18 ;
    END
  END Y
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.745 2.58 1.61 2.58 1.61 2.61 1.31 2.61 1.31 2.275 1.13 2.275 1.13 2.215 1.16 2.215 1.16 1.93 0.81 1.93 0.81 2.265 0.75 2.265 0.75 1.87 1.22 1.87 1.22 2.215 1.37 2.215 1.37 2.49 1.61 2.49 1.61 2.52 1.685 2.52 1.685 1.95 1.745 1.95 ;
    END
  END ExtVDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.57 2.455 0.81 2.575 ;
    END
  END A
  PIN ISOn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.29629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.78 2.66 1 2.78 ;
    END
  END ISOn
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 3.48 0 3.48 0 3.36 1.045 3.36 1.045 3.005 1.105 3.005 1.105 3.36 1.685 3.36 1.685 2.92 1.745 2.92 1.745 3.36 2.8 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 2.8 0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 2.8 1.77 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.83 2.79 1.14 2.79 1.14 2.935 0.795 2.935 0.795 3.15 0.735 3.15 0.735 2.875 1.08 2.875 1.08 2.425 0.955 2.425 0.955 2.05 1.015 2.05 1.015 2.365 1.14 2.365 1.14 2.73 1.83 2.73 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END ISONLX1_OFF

MACRO ISONLX1_ON
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ISONLX1_ON 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.522 LAYER Metal1 ;
    ANTENNADIFFAREA 0.6139 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 17.84615375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 149.64102575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.165 1.11 1.055 1.11 1.055 1.465 0.995 1.465 0.995 0.245 1.055 0.245 1.055 0.975 1.165 0.975 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.14 1.65 0.14 1.25 0.2 1.25 0.2 1.65 0.55 1.65 0.55 1.25 0.61 1.25 0.61 1.65 0.79 1.65 0.79 1.075 0.85 1.075 0.85 1.65 1.2 1.65 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.68518525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.505 0.79 0.765 0.945 ;
    END
  END A
  PIN ISOn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.035 0.6 0.25 0.75 ;
    END
  END ISOn
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.85 0.06 0.85 0.505 0.79 0.505 0.79 0.06 0.3 0.06 0.3 0.39 0.24 0.39 0.24 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.935 0.68 0.405 0.68 0.405 1.465 0.345 1.465 0.345 0.62 0.55 0.62 0.55 0.245 0.61 0.245 0.61 0.62 0.935 0.62 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END ISONLX1_ON

MACRO LSHL_ISOH_X1_FROM_OFF
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSHL_ISOH_X1_FROM_OFF 0 0 ;
  SIZE 2.8 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.745 2.39 1.685 2.39 1.685 1.93 1.095 1.93 1.095 2.49 1.24 2.49 1.24 2.63 0.835 2.63 0.835 2.49 1.035 2.49 1.035 1.87 1.745 1.87 ;
    END
  END ExtVDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.83333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 2.485 0.765 2.63 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9839 LAYER Metal1 ;
    ANTENNADIFFAREA 0.9138 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0702 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.0156695 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 113.5470085 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.97 3.01 1.95 3.01 1.95 3.14 1.89 3.14 1.89 3.01 1.84 3.01 1.84 2.88 1.89 2.88 1.89 2.51 1.48 2.51 1.48 2 1.54 2 1.54 2.45 1.89 2.45 1.89 2 1.95 2 1.95 2.88 1.97 2.88 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 3.48 0 3.48 0 3.36 0.145 3.36 0.145 2.88 0.205 2.88 0.205 3.36 1.24 3.36 1.24 3.02 1.3 3.02 1.3 3.36 2.8 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 2.8 0.06 ;
    END
  END VSS
  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.18 2.295 0.365 2.44 ;
    END
  END ISO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 2.8 1.77 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.815 2.68 1.395 2.68 1.395 2.795 0.65 2.795 0.65 3.025 0.59 3.025 0.59 2.735 1.335 2.735 1.335 2.245 1.24 2.245 1.24 2 1.3 2 1.3 2.185 1.395 2.185 1.395 2.62 1.815 2.62 ;
      POLYGON 1.745 3.14 1.445 3.14 1.445 2.95 1.095 2.95 1.095 3.14 1.005 3.14 1.005 3.03 0.855 3.03 0.855 3.025 0.795 3.025 0.795 2.88 1.745 2.88 ;
      POLYGON 1.055 3.275 0.86 3.275 0.86 3.195 0.35 3.195 0.35 2.83 0.425 2.83 0.425 2.26 0.83 2.26 0.83 2 0.89 2 0.89 2.32 0.485 2.32 0.485 2.89 0.41 2.89 0.41 3.135 0.92 3.135 0.92 3.215 1.055 3.215 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSHL_ISOH_X1_FROM_OFF

MACRO LSHL_ISOH_X1_TO_ON
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSHL_ISOH_X1_TO_ON 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 0.79 0.765 0.93 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2371 LAYER Metal1 ;
    ANTENNADIFFAREA 1.0626 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0702 LAYER Metal1 ;
      ANTENNAMAXAREACAR 17.622507 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 127.30769225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.965 1.3 1.95 1.3 1.95 1.42 1.89 1.42 1.89 1.3 1.835 1.3 1.835 0.885 1.54 0.885 1.54 1.42 1.48 1.42 1.48 0.825 1.835 0.825 1.835 0.79 1.89 0.79 1.89 0.28 1.95 0.28 1.95 0.79 1.965 0.79 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 1.3 0.06 1.3 0.4 1.24 0.4 1.24 0.06 0.205 0.06 0.205 0.54 0.145 0.54 0.145 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
  END VSS
  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.9444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.135 0.98 0.365 1.125 ;
    END
  END ISO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 1.035 1.65 1.035 1.205 1.095 1.205 1.095 1.65 1.685 1.65 1.685 1.03 1.745 1.03 1.745 1.65 2.2 1.65 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.82 0.695 1.395 0.695 1.395 1.235 1.3 1.235 1.3 1.42 1.24 1.42 1.24 1.175 1.335 1.175 1.335 0.67 0.59 0.67 0.59 0.395 0.65 0.395 0.65 0.61 1.395 0.61 1.395 0.635 1.82 0.635 ;
      POLYGON 1.745 0.54 0.795 0.54 0.795 0.395 0.855 0.395 0.855 0.39 1.005 0.39 1.005 0.28 1.095 0.28 1.095 0.47 1.445 0.47 1.445 0.28 1.745 0.28 ;
      POLYGON 1.055 0.205 0.92 0.205 0.92 0.285 0.41 0.285 0.41 0.48 0.515 0.48 0.515 1.1 0.89 1.1 0.89 1.42 0.83 1.42 0.83 1.16 0.455 1.16 0.455 0.54 0.35 0.54 0.35 0.225 0.86 0.225 0.86 0.145 1.055 0.145 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSHL_ISOH_X1_TO_ON

MACRO LSHL_ISOL_X1_FROM_OFF
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSHL_ISOL_X1_FROM_OFF 0 0 ;
  SIZE 2.8 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.745 2.39 1.685 2.39 1.685 1.93 1.095 1.93 1.095 2.5 1.24 2.5 1.24 2.63 0.835 2.63 0.835 2.5 1.035 2.5 1.035 1.87 1.745 1.87 ;
    END
  END ExtVDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.29629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 2.31 0.765 2.48 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.98735 LAYER Metal1 ;
    ANTENNADIFFAREA 0.89225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.062325 LAYER Metal1 ;
      ANTENNAMAXAREACAR 15.8419575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 127.2683515 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.965 2.82 1.95 2.82 1.95 3.14 1.89 3.14 1.89 2.82 1.835 2.82 1.835 2.69 1.89 2.69 1.89 2 1.95 2 1.95 2.69 1.965 2.69 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 3.48 0 3.48 0 3.36 0.145 3.36 0.145 2.88 0.205 2.88 0.205 3.36 1.24 3.36 1.24 3.02 1.3 3.02 1.3 3.36 1.685 3.36 1.685 2.88 1.745 2.88 1.745 3.36 2.8 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 2.8 0.06 ;
    END
  END VSS
  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.64814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 2.105 0.365 2.25 ;
    END
  END ISO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 2.8 1.77 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.82 2.58 1.395 2.58 1.395 2.79 0.65 2.79 0.65 3.025 0.59 3.025 0.59 2.73 1.335 2.73 1.335 2.215 1.24 2.215 1.24 2 1.3 2 1.3 1.995 1.45 1.995 1.45 2 1.51 2 1.51 2.215 1.395 2.215 1.395 2.52 1.82 2.52 ;
      POLYGON 1.505 3.14 1.445 3.14 1.445 2.95 1.095 2.95 1.095 3.14 1.005 3.14 1.005 3.03 0.855 3.03 0.855 3.025 0.795 3.025 0.795 2.88 1.505 2.88 ;
      POLYGON 1.055 3.275 0.86 3.275 0.86 3.195 0.35 3.195 0.35 2.88 0.425 2.88 0.425 2.155 0.83 2.155 0.83 2 0.89 2 0.89 2.215 0.485 2.215 0.485 2.94 0.41 2.94 0.41 3.135 0.92 3.135 0.92 3.215 1.055 3.215 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSHL_ISOL_X1_FROM_OFF

MACRO LSHL_ISOL_X1_TO_ON
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSHL_ISOL_X1_TO_ON 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 0.79 0.765 0.93 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0862 LAYER Metal1 ;
    ANTENNADIFFAREA 1.07115 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.062325 LAYER Metal1 ;
      ANTENNAMAXAREACAR 17.4279985 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 132.17809875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.965 1.11 1.95 1.11 1.95 1.42 1.89 1.42 1.89 1.11 1.835 1.11 1.835 0.79 1.89 0.79 1.89 0.28 1.95 0.28 1.95 0.79 1.965 0.79 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 1.745 0.06 1.745 0.54 1.685 0.54 1.685 0.06 1.3 0.06 1.3 0.4 1.24 0.4 1.24 0.06 0.205 0.06 0.205 0.54 0.145 0.54 0.145 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
  END VSS
  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.205 0.6 0.365 0.765 ;
    END
  END ISO
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 1.035 1.65 1.035 1.205 1.095 1.205 1.095 1.65 1.685 1.65 1.685 1.03 1.745 1.03 1.745 1.65 2.2 1.65 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.82 0.71 1.395 0.71 1.395 1.205 1.51 1.205 1.51 1.42 1.45 1.42 1.45 1.425 1.3 1.425 1.3 1.42 1.24 1.42 1.24 1.205 1.335 1.205 1.335 0.71 0.59 0.71 0.59 0.395 0.65 0.395 0.65 0.65 1.82 0.65 ;
      POLYGON 1.505 0.54 0.795 0.54 0.795 0.395 0.855 0.395 0.855 0.39 1.005 0.39 1.005 0.28 1.095 0.28 1.095 0.47 1.445 0.47 1.445 0.28 1.505 0.28 ;
      POLYGON 1.055 0.205 0.92 0.205 0.92 0.285 0.41 0.285 0.41 0.48 0.485 0.48 0.485 1.1 0.89 1.1 0.89 1.42 0.83 1.42 0.83 1.16 0.425 1.16 0.425 0.54 0.35 0.54 0.35 0.225 0.86 0.225 0.86 0.145 1.055 0.145 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSHL_ISOL_X1_TO_ON

MACRO LSHL_ISONH_X1_FROM_OFF
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSHL_ISONH_X1_FROM_OFF 0 0 ;
  SIZE 2.8 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.745 2.39 1.685 2.39 1.685 1.93 1.095 1.93 1.095 2.49 1.24 2.49 1.24 2.61 0.88 2.61 0.88 2.49 1.035 2.49 1.035 1.87 1.745 1.87 ;
    END
  END ExtVDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.27777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 2.485 0.74 2.625 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7979 LAYER Metal1 ;
    ANTENNADIFFAREA 0.8388 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 27.2786325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 210.923077 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.95 3.185 1.89 3.185 1.89 2.53 1.48 2.53 1.48 2 1.54 2 1.54 2.47 1.89 2.47 1.89 2 1.95 2 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 3.48 0 3.48 0 3.36 1.24 3.36 1.24 3.065 1.3 3.065 1.3 3.36 2.8 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 2.8 0.06 ;
    END
  END VSS
  PIN ISOn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04095 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.34432225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.505 2.59 1.725 2.69 ;
    END
  END ISOn
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 2.8 1.77 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.82 2.845 0.65 2.845 0.65 3.07 0.59 3.07 0.59 2.785 1.335 2.785 1.335 2.245 1.24 2.245 1.24 2 1.3 2 1.3 2.185 1.395 2.185 1.395 2.785 1.82 2.785 ;
      POLYGON 1.745 3.185 1.445 3.185 1.445 2.995 1.095 2.995 1.095 3.185 1.005 3.185 1.005 3.075 0.855 3.075 0.855 3.07 0.795 3.07 0.795 2.925 1.745 2.925 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSHL_ISONH_X1_FROM_OFF

MACRO LSHL_ISONH_X1_TO_ON
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSHL_ISONH_X1_TO_ON 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.83333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.145 1.005 0.36 1.105 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8108 LAYER Metal1 ;
    ANTENNADIFFAREA 0.8916 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 27.719658 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 205.84615375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.59 1.42 1.53 1.42 1.53 0.95 1.18 0.95 1.18 1.42 1.12 1.42 1.12 0.89 1.53 0.89 1.53 0.28 1.59 0.28 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 0.94 0.06 0.94 0.4 0.88 0.4 0.88 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
  END VSS
  PIN ISOn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04095 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.4175825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.6 0.83 0.83 0.93 ;
    END
  END ISOn
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.675 1.65 0.675 1.205 0.735 1.205 0.735 1.65 1.325 1.65 1.325 1.03 1.385 1.03 1.385 1.65 1.8 1.65 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.46 0.71 1.035 0.71 1.035 1.235 0.94 1.235 0.94 1.42 0.88 1.42 0.88 1.175 0.975 1.175 0.975 0.71 0.23 0.71 0.23 0.395 0.29 0.395 0.29 0.65 1.46 0.65 ;
      POLYGON 1.385 0.54 0.435 0.54 0.435 0.395 0.495 0.395 0.495 0.39 0.645 0.39 0.645 0.28 0.735 0.28 0.735 0.47 1.085 0.47 1.085 0.28 1.385 0.28 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSHL_ISONH_X1_TO_ON

MACRO LSHL_ISONL_X1_FROM_OFF
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSHL_ISONL_X1_FROM_OFF 0 0 ;
  SIZE 2.8 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.745 2.39 1.685 2.39 1.685 1.93 1.095 1.93 1.095 2.49 1.24 2.49 1.24 2.61 0.88 2.61 0.88 2.49 1.035 2.49 1.035 1.87 1.745 1.87 ;
    END
  END ExtVDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.27777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.595 2.485 0.74 2.625 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8045 LAYER Metal1 ;
    ANTENNADIFFAREA 0.81725 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 27.5042735 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 208.82051275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.89 2 1.95 3.14 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 3.48 0 3.48 0 3.36 1.24 3.36 1.24 3.02 1.3 3.02 1.3 3.36 1.685 3.36 1.685 2.88 1.745 2.88 1.745 3.36 2.8 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 2.8 0.06 ;
    END
  END VSS
  PIN ISOn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.033075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.675737 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.48 2.49 1.655 2.61 ;
    END
  END ISOn
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 2.8 1.77 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.82 2.77 0.65 2.77 0.65 3.025 0.59 3.025 0.59 2.71 1.335 2.71 1.335 2.215 1.24 2.215 1.24 2 1.3 2 1.3 1.995 1.45 1.995 1.45 2 1.51 2 1.51 2.215 1.395 2.215 1.395 2.71 1.82 2.71 ;
      POLYGON 1.505 3.14 1.445 3.14 1.445 2.95 1.095 2.95 1.095 3.14 1.005 3.14 1.005 3.03 0.855 3.03 0.855 3.025 0.795 3.025 0.795 2.88 1.505 2.88 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSHL_ISONL_X1_FROM_OFF

MACRO LSHL_ISONL_X1_TO_ON
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSHL_ISONL_X1_TO_ON 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.27777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.175 0.795 0.32 0.935 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8174 LAYER Metal1 ;
    ANTENNADIFFAREA 0.87005 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 27.94529925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 204.20512825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.47 0.28 1.53 1.42 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.325 0.06 1.325 0.54 1.265 0.54 1.265 0.06 0.88 0.06 0.88 0.4 0.82 0.4 0.82 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
  END VSS
  PIN ISOn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.033075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.537415 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.87 0.925 0.97 ;
    END
  END ISOn
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.615 1.65 0.615 1.205 0.675 1.205 0.675 1.65 1.265 1.65 1.265 1.03 1.325 1.03 1.325 1.65 1.8 1.65 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.4 0.71 1.09 0.71 1.09 1.42 1.03 1.42 1.03 1.425 0.88 1.425 0.88 1.42 0.82 1.42 0.82 1.205 1.03 1.205 1.03 0.71 0.17 0.71 0.17 0.395 0.23 0.395 0.23 0.65 1.4 0.65 ;
      POLYGON 1.085 0.54 0.375 0.54 0.375 0.395 0.435 0.395 0.435 0.39 0.585 0.39 0.585 0.28 0.675 0.28 0.675 0.47 1.025 0.47 1.025 0.28 1.085 0.28 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSHL_ISONL_X1_TO_ON

MACRO LSHLX1_FROM
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSHLX1_FROM 0 0 ;
  SIZE 2.6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.575 2.585 1.365 2.585 1.365 2.63 0.955 2.63 0.955 2.035 1.015 2.035 1.015 2.49 1.365 2.49 1.365 2.525 1.515 2.525 1.515 2.055 1.575 2.055 ;
    END
  END ExtVDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.4814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.37 2.31 0.59 2.44 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6028 LAYER Metal1 ;
    ANTENNADIFFAREA 0.638 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 20.608547 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 161.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.965 2.82 1.78 2.82 1.78 3.16 1.72 3.16 1.72 2.055 1.78 2.055 1.78 2.69 1.965 2.69 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 3.48 0 3.48 0 3.36 0.955 3.36 0.955 2.97 1.015 2.97 1.015 3.36 1.515 3.36 1.515 2.9 1.575 2.9 1.575 3.36 2.6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 2.6 0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 2.6 1.77 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.635 2.795 0.81 2.795 0.81 3.115 0.75 3.115 0.75 2.035 0.81 2.035 0.81 2.735 1.635 2.735 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSHLX1_FROM

MACRO LSHLX1_TO
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSHLX1_TO 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.77 0 1.77 0 1.65 0.375 1.65 0.375 1.03 0.435 1.03 0.435 1.65 0.8 1.65 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.388889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.79 0.45 0.92 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3456 LAYER Metal1 ;
    ANTENNADIFFAREA 0.4424 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.8153845 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 103.12820525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.765 0.73 0.64 0.73 0.64 1.42 0.58 1.42 0.58 0.27 0.64 0.27 0.64 0.6 0.765 0.6 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 0.06 0.435 0.06 0.435 0.53 0.375 0.53 0.375 0.06 0 0.06 0 -0.06 0.8 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.495 0.675 0.175 0.675 0.175 1.12 0.2 1.12 0.2 1.335 0.115 1.335 0.115 0.335 0.2 0.335 0.2 0.48 0.175 0.48 0.175 0.615 0.495 0.615 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSHLX1_TO

MACRO LSLH_ISOH_X1_FROM_OFF
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSLH_ISOH_X1_FROM_OFF 0 0 ;
  SIZE 4 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 0.295 1.77 0.295 2.255 0.235 2.255 0.235 1.77 0 1.77 0 1.65 4 1.65 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0513 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.6959065 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.22 2.675 0.365 2.82 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6379 LAYER Metal1 ;
    ANTENNADIFFAREA 1.6996 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.14805 LAYER Metal1 ;
      ANTENNAMAXAREACAR 17.81762925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 145.5116515 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.365 2.25 3.235 2.25 3.235 3.185 3.175 3.185 3.175 1.95 2.845 1.95 2.845 1.89 3.365 1.89 ;
    END
  END Y
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.03 2.46 2.97 2.46 2.97 2.265 2.59 2.265 2.59 2.49 2.765 2.49 2.765 2.63 2.435 2.63 2.435 2.5 2.465 2.5 2.465 2.49 2.53 2.49 2.53 2.265 2.27 2.265 2.27 1.93 1.45 1.93 1.45 2.265 1.39 2.265 1.39 1.87 2.33 1.87 2.33 2.205 2.53 2.205 2.53 2 2.59 2 2.59 2.205 2.97 2.205 2.97 2.07 3.03 2.07 ;
    END
  END ExtVDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.36 4 3.48 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.015 0.06 3.015 0.51 2.955 0.51 2.955 0.06 2.605 0.06 2.605 0.51 2.545 0.51 2.545 0.06 2.195 0.06 2.195 0.51 2.135 0.51 2.135 0.06 1.5 0.06 1.5 0.415 1.44 0.415 1.44 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
  END VSS
  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.235 0.6 1.565 0.73 ;
    END
  END ISO
  OBS
    LAYER Metal1 ;
      POLYGON 3.09 2.76 3.06 2.76 3.06 2.79 2.635 2.79 2.635 3.13 2.575 3.13 2.575 2.79 2.225 2.79 2.225 3.13 2.165 3.13 2.165 2.53 1.595 2.53 1.595 2.05 1.655 2.05 1.655 2.47 2.265 2.47 2.265 2.53 2.225 2.53 2.225 2.73 2.97 2.73 2.97 2.7 3.09 2.7 ;
      POLYGON 3.03 3.255 0.235 3.255 0.235 2.98 0.295 2.98 0.295 3.195 0.93 3.195 0.93 1.97 0.99 1.97 0.99 3.195 1.55 3.195 1.55 2.87 1.61 2.87 1.61 3.195 1.96 3.195 1.96 2.87 2.02 2.87 2.02 3.195 2.37 3.195 2.37 2.87 2.43 2.87 2.43 3.195 2.97 3.195 2.97 2.925 3.03 2.925 ;
      POLYGON 2.96 1.555 2.79 1.555 2.79 0.955 2.85 0.955 2.85 1.495 2.96 1.495 ;
      POLYGON 2.81 0.855 2.4 0.855 2.4 0.915 0.99 0.915 0.99 1.515 0.93 1.515 0.93 0.855 2.34 0.855 2.34 0.25 2.4 0.25 2.4 0.795 2.75 0.795 2.75 0.25 2.81 0.25 ;
      POLYGON 2.645 1.53 1.44 1.53 1.44 1.13 1.5 1.13 1.5 1.47 2.585 1.47 2.585 0.955 2.645 0.955 ;
      POLYGON 2.125 2.39 1.81 2.39 1.81 2.33 2.065 2.33 2.065 2.05 2.125 2.05 ;
      POLYGON 2.08 1.035 1.705 1.035 1.705 1.345 1.645 1.345 1.645 0.975 2.08 0.975 ;
      POLYGON 1.91 0.64 1.645 0.64 1.645 0.27 1.705 0.27 1.705 0.58 1.91 0.58 ;
      POLYGON 1.815 3.13 1.755 3.13 1.755 2.74 1.405 2.74 1.405 3.13 1.345 3.13 1.345 2.335 1.405 2.335 1.405 2.68 1.815 2.68 ;
      POLYGON 0.62 2.855 0.5 2.855 0.5 3.125 0.44 3.125 0.44 2.04 0.5 2.04 0.5 2.795 0.62 2.795 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSLH_ISOH_X1_FROM_OFF

MACRO LSLH_ISOH_X1_TO_ON
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSLH_ISOH_X1_TO_ON 0 0 ;
  SIZE 4 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 2.93 1.77 2.93 2.175 3.57 2.175 3.57 2.09 3.63 2.09 3.63 2.48 3.57 2.48 3.57 2.235 2.87 2.235 2.87 1.77 2.05 1.77 2.05 2.205 1.99 2.205 1.99 1.77 0 1.77 0 1.65 2.345 1.65 2.345 1.185 2.405 1.185 2.405 1.65 3.195 1.65 3.195 0.96 3.255 0.96 3.255 1.65 4 1.65 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0513 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.04678375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.62 2.71 0.85 2.83 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4696 LAYER Metal1 ;
    ANTENNADIFFAREA 1.68655 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.14805 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.680851 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 136.98074975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.835 3.04 3.775 3.04 3.775 1.955 3.37 1.955 3.37 1.895 3.835 1.895 ;
    END
  END Y
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.085 2.61 0.785 2.61 0.785 2.49 0.835 2.49 0.835 1.975 0.895 1.975 0.895 2.49 1.085 2.49 ;
    END
  END ExtVDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.36 4 3.48 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.46 0.06 3.46 0.535 3.4 0.535 3.4 0.06 3.05 0.06 3.05 0.535 2.99 0.535 2.99 0.06 2.64 0.06 2.64 0.535 2.58 0.535 2.58 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
  END VSS
  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.5555555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.275 0.965 2.455 1.085 ;
    END
  END ISO
  OBS
    LAYER Metal1 ;
      POLYGON 3.7 2.66 3.235 2.66 3.235 3.04 3.175 3.04 3.175 2.66 2.825 2.66 2.825 3.04 2.765 3.04 2.765 2.45 2.195 2.45 2.195 1.99 2.255 1.99 2.255 2.39 2.705 2.39 2.705 2.37 2.825 2.37 2.825 2.6 3.7 2.6 ;
      POLYGON 3.63 3.245 0.835 3.245 0.835 2.95 0.895 2.95 0.895 3.185 1.685 3.185 1.685 1.925 1.745 1.925 1.745 3.185 2.15 3.185 2.15 2.78 2.21 2.78 2.21 3.185 2.56 3.185 2.56 2.78 2.62 2.78 2.62 3.185 2.97 3.185 2.97 2.78 3.03 2.78 3.03 3.185 3.57 3.185 3.57 2.78 3.63 2.78 ;
      POLYGON 3.525 1.57 3.4 1.57 3.4 0.96 3.46 0.96 3.46 1.51 3.525 1.51 ;
      POLYGON 3.255 0.87 1.745 0.87 1.745 1.465 1.685 1.465 1.685 0.81 2.785 0.81 2.785 0.275 2.845 0.275 2.845 0.81 3.195 0.81 3.195 0.275 3.255 0.275 ;
      POLYGON 2.77 1.085 2.61 1.085 2.61 1.4 2.55 1.4 2.55 1.025 2.77 1.025 ;
      POLYGON 2.725 2.21 2.41 2.21 2.41 2.15 2.665 2.15 2.665 1.99 2.725 1.99 ;
      POLYGON 2.715 0.695 2.345 0.695 2.345 0.32 2.405 0.32 2.405 0.635 2.715 0.635 ;
      POLYGON 2.415 3.04 2.355 3.04 2.355 2.66 2.005 2.66 2.005 3.04 1.945 3.04 1.945 2.275 2.005 2.275 2.005 2.6 2.415 2.6 ;
      POLYGON 1.57 2.74 1.51 2.74 1.51 3.01 1.1 3.01 1.1 3.095 1.04 3.095 1.04 2.95 1.45 2.95 1.45 2.19 1.04 2.19 1.04 1.975 1.1 1.975 1.1 2.13 1.51 2.13 1.51 2.68 1.57 2.68 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSLH_ISOH_X1_TO_ON

MACRO LSLH_ISOL_X1_FROM_OFF
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSLH_ISOL_X1_FROM_OFF 0 0 ;
  SIZE 4 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 0.295 1.77 0.295 2.255 0.235 2.255 0.235 1.77 0 1.77 0 1.65 4 1.65 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0513 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.6959065 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.22 2.675 0.365 2.82 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.06665 LAYER Metal1 ;
    ANTENNADIFFAREA 2.1306 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.140175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 21.87729625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 167.8758695 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.365 2.44 3.235 2.44 3.235 3.185 3.175 3.185 3.175 1.955 3.235 1.955 3.235 2.105 3.365 2.105 ;
    END
  END Y
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.03 2.345 2.97 2.345 2.97 2.265 2.645 2.265 2.645 2.49 2.765 2.49 2.765 2.63 2.435 2.63 2.435 2.49 2.585 2.49 2.585 2.265 2.27 2.265 2.27 1.93 1.45 1.93 1.45 2.265 1.39 2.265 1.39 1.87 2.33 1.87 2.33 2.205 2.585 2.205 2.585 2 2.645 2 2.645 2.205 2.97 2.205 2.97 1.955 3.03 1.955 ;
    END
  END ExtVDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 3.48 0 3.48 0 3.36 2.97 3.36 2.97 2.925 3.03 2.925 3.03 3.36 4 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.015 0.06 3.015 0.51 2.955 0.51 2.955 0.06 2.605 0.06 2.605 0.51 2.545 0.51 2.545 0.06 2.195 0.06 2.195 0.51 2.135 0.51 2.135 0.06 1.5 0.06 1.5 0.415 1.44 0.415 1.44 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
  END VSS
  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.185 0.55 1.565 0.73 ;
    END
  END ISO
  OBS
    LAYER Metal1 ;
      POLYGON 3.165 1.545 2.79 1.545 2.79 1.055 2.85 1.055 2.85 1.485 3.165 1.485 ;
      POLYGON 3.09 2.76 3.06 2.76 3.06 2.79 2.635 2.79 2.635 3.13 2.575 3.13 2.575 2.79 2.225 2.79 2.225 3.13 2.165 3.13 2.165 2.53 1.595 2.53 1.595 2.05 1.655 2.05 1.655 2.47 2.265 2.47 2.265 2.53 2.225 2.53 2.225 2.73 2.97 2.73 2.97 2.7 3.09 2.7 ;
      POLYGON 2.81 0.84 2.4 0.84 2.4 0.915 0.99 0.915 0.99 1.515 0.93 1.515 0.93 0.855 2.34 0.855 2.34 0.25 2.4 0.25 2.4 0.78 2.75 0.78 2.75 0.25 2.81 0.25 ;
      POLYGON 2.645 1.575 2.585 1.575 2.585 1.53 1.44 1.53 1.44 1.13 1.5 1.13 1.5 1.47 2.585 1.47 2.585 1.055 2.645 1.055 ;
      POLYGON 2.43 3.255 0.235 3.255 0.235 2.98 0.295 2.98 0.295 3.195 0.93 3.195 0.93 1.97 0.99 1.97 0.99 3.195 1.55 3.195 1.55 2.87 1.61 2.87 1.61 3.195 1.96 3.195 1.96 2.87 2.02 2.87 2.02 3.195 2.37 3.195 2.37 2.87 2.43 2.87 ;
      POLYGON 2.125 2.39 1.81 2.39 1.81 2.33 2.065 2.33 2.065 2.05 2.125 2.05 ;
      POLYGON 2.08 1.035 1.705 1.035 1.705 1.345 1.645 1.345 1.645 0.975 2.08 0.975 ;
      POLYGON 1.91 0.64 1.705 0.64 1.705 0.415 1.645 0.415 1.645 0.27 1.705 0.27 1.705 0.355 1.765 0.355 1.765 0.58 1.91 0.58 ;
      POLYGON 1.815 3.13 1.755 3.13 1.755 2.74 1.405 2.74 1.405 3.13 1.345 3.13 1.345 2.335 1.405 2.335 1.405 2.68 1.815 2.68 ;
      POLYGON 0.62 2.85 0.5 2.85 0.5 3.125 0.44 3.125 0.44 2.04 0.5 2.04 0.5 2.79 0.62 2.79 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSLH_ISOL_X1_FROM_OFF

MACRO LSLH_ISOL_X1_TO_ON
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSLH_ISOL_X1_TO_ON 0 0 ;
  SIZE 4 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 3.555 1.77 3.555 2.37 3.495 2.37 3.495 1.77 2.93 1.77 2.93 2.205 2.87 2.205 2.87 1.77 2.05 1.77 2.05 2.205 1.99 2.205 1.99 1.77 0 1.77 0 1.65 2.345 1.65 2.345 1.185 2.405 1.185 2.405 1.65 3.195 1.65 3.195 1.135 3.255 1.135 3.255 1.65 4 1.65 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0513 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.0760235 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 2.69 0.85 2.83 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9032 LAYER Metal1 ;
    ANTENNADIFFAREA 2.11755 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.140175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 20.71125375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 155.848047 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.81 2.44 3.76 2.44 3.76 3.04 3.7 3.04 3.7 2.44 3.63 2.44 3.63 2.105 3.7 2.105 3.7 1.98 3.76 1.98 3.76 2.105 3.81 2.105 ;
    END
  END Y
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.165 2.63 0.785 2.63 0.785 2.49 0.835 2.49 0.835 1.975 0.895 1.975 0.895 2.49 1.165 2.49 ;
    END
  END ExtVDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 3.48 0 3.48 0 3.36 3.495 3.36 3.495 2.78 3.555 2.78 3.555 3.36 4 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.46 0.06 3.46 0.535 3.4 0.535 3.4 0.06 3.05 0.06 3.05 0.535 2.99 0.535 2.99 0.06 2.64 0.06 2.64 0.535 2.58 0.535 2.58 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
  END VSS
  PIN ISO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.5555555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.275 0.965 2.455 1.085 ;
    END
  END ISO
  OBS
    LAYER Metal1 ;
      POLYGON 3.69 1.475 3.4 1.475 3.4 1.135 3.46 1.135 3.46 1.415 3.69 1.415 ;
      POLYGON 3.625 2.66 3.235 2.66 3.235 3.04 3.175 3.04 3.175 2.66 2.825 2.66 2.825 3.04 2.765 3.04 2.765 2.45 2.195 2.45 2.195 1.99 2.255 1.99 2.255 2.39 2.705 2.39 2.705 2.37 2.825 2.37 2.825 2.6 3.625 2.6 ;
      POLYGON 3.255 0.87 1.745 0.87 1.745 1.465 1.685 1.465 1.685 0.81 2.785 0.81 2.785 0.275 2.845 0.275 2.845 0.81 3.195 0.81 3.195 0.275 3.255 0.275 ;
      POLYGON 3.03 3.245 0.835 3.245 0.835 2.95 0.895 2.95 0.895 3.185 1.685 3.185 1.685 1.925 1.745 1.925 1.745 3.185 2.15 3.185 2.15 2.78 2.21 2.78 2.21 3.185 2.56 3.185 2.56 2.78 2.62 2.78 2.62 3.185 2.97 3.185 2.97 2.78 3.03 2.78 ;
      POLYGON 2.77 1.085 2.61 1.085 2.61 1.4 2.55 1.4 2.55 1.025 2.77 1.025 ;
      POLYGON 2.725 2.21 2.41 2.21 2.41 2.15 2.665 2.15 2.665 1.99 2.725 1.99 ;
      POLYGON 2.715 0.695 2.345 0.695 2.345 0.32 2.405 0.32 2.405 0.635 2.715 0.635 ;
      POLYGON 2.415 3.04 2.355 3.04 2.355 2.66 2.005 2.66 2.005 3.04 1.945 3.04 1.945 2.275 2.005 2.275 2.005 2.6 2.415 2.6 ;
      POLYGON 1.57 2.74 1.51 2.74 1.51 3.01 1.1 3.01 1.1 3.095 1.04 3.095 1.04 2.95 1.45 2.95 1.45 2.19 1.04 2.19 1.04 1.975 1.1 1.975 1.1 2.13 1.51 2.13 1.51 2.68 1.57 2.68 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSLH_ISOL_X1_TO_ON

MACRO LSLH_ISONH_X1_FROM_OFF
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSLH_ISONH_X1_FROM_OFF 0 0 ;
  SIZE 4 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 0.295 1.77 0.295 2.255 0.235 2.255 0.235 1.77 0 1.77 0 1.65 4 1.65 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0513 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.72514625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.22 2.67 0.365 2.82 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4542 LAYER Metal1 ;
    ANTENNADIFFAREA 1.5988 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0837 LAYER Metal1 ;
      ANTENNAMAXAREACAR 29.321386 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 234.014337 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.375 2.455 3.235 2.455 3.235 3.185 3.175 3.185 3.175 1.935 2.765 1.935 2.765 1.875 3.235 1.875 3.235 2.085 3.375 2.085 ;
    END
  END Y
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.03 2.41 2.97 2.41 2.97 2.265 2.645 2.265 2.645 2.49 2.765 2.49 2.765 2.63 2.435 2.63 2.435 2.49 2.585 2.49 2.585 2.265 2.27 2.265 2.27 1.93 1.45 1.93 1.45 2.265 1.39 2.265 1.39 1.87 2.33 1.87 2.33 2.205 2.585 2.205 2.585 2 2.645 2 2.645 2.205 2.97 2.205 2.97 2.02 3.03 2.02 ;
    END
  END ExtVDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.36 4 3.48 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.015 0.06 3.015 0.51 2.955 0.51 2.955 0.06 2.605 0.06 2.605 0.51 2.545 0.51 2.545 0.06 2.195 0.06 2.195 0.51 2.135 0.51 2.135 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
  END VSS
  PIN ISOn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06435 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.63170175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.01 0.73 3.26 0.83 ;
    END
  END ISOn
  OBS
    LAYER Metal1 ;
      POLYGON 3.09 2.76 3.06 2.76 3.06 2.79 2.635 2.79 2.635 3.13 2.575 3.13 2.575 2.79 2.225 2.79 2.225 3.13 2.165 3.13 2.165 2.53 1.595 2.53 1.595 2.05 1.655 2.05 1.655 2.47 2.265 2.47 2.265 2.53 2.225 2.53 2.225 2.73 2.97 2.73 2.97 2.7 3.09 2.7 ;
      POLYGON 3.03 3.255 0.235 3.255 0.235 2.98 0.295 2.98 0.295 3.195 0.93 3.195 0.93 1.97 0.99 1.97 0.99 3.195 1.55 3.195 1.55 2.87 1.61 2.87 1.61 3.195 1.96 3.195 1.96 2.87 2.02 2.87 2.02 3.195 2.37 3.195 2.37 2.87 2.43 2.87 2.43 3.195 2.97 3.195 2.97 2.925 3.03 2.925 ;
      RECT 2.79 0.905 2.85 1.57 ;
      POLYGON 2.81 0.72 0.99 0.72 0.99 1.515 0.93 1.515 0.93 0.66 2.34 0.66 2.34 0.25 2.4 0.25 2.4 0.66 2.75 0.66 2.75 0.25 2.81 0.25 ;
      RECT 2.585 0.905 2.645 1.575 ;
      POLYGON 2.125 2.39 1.81 2.39 1.81 2.33 2.065 2.33 2.065 2.05 2.125 2.05 ;
      POLYGON 1.815 3.13 1.755 3.13 1.755 2.74 1.405 2.74 1.405 3.13 1.345 3.13 1.345 2.335 1.405 2.335 1.405 2.68 1.815 2.68 ;
      POLYGON 0.62 2.855 0.5 2.855 0.5 3.125 0.44 3.125 0.44 2.04 0.5 2.04 0.5 2.795 0.62 2.795 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSLH_ISONH_X1_FROM_OFF

MACRO LSLH_ISONH_X1_TO_ON
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSLH_ISONH_X1_TO_ON 0 0 ;
  SIZE 4 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 2.935 1.77 2.935 2.175 3.575 2.175 3.575 2.09 3.635 2.09 3.635 2.48 3.575 2.48 3.575 2.235 2.875 2.235 2.875 1.77 2.055 1.77 2.055 2.205 1.995 2.205 1.995 1.77 0 1.77 0 1.65 3.2 1.65 3.2 0.96 3.26 0.96 3.26 1.65 4 1.65 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0513 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.04678375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.625 2.71 0.855 2.83 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3586 LAYER Metal1 ;
    ANTENNADIFFAREA 1.5988 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0837 LAYER Metal1 ;
      ANTENNAMAXAREACAR 28.1792115 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 228.172043 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.84 3.04 3.78 3.04 3.78 1.955 3.375 1.955 3.375 1.895 3.84 1.895 ;
    END
  END Y
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.09 2.61 0.79 2.61 0.79 2.49 0.84 2.49 0.84 1.975 0.9 1.975 0.9 2.49 1.09 2.49 ;
    END
  END ExtVDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 3.36 4 3.48 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.465 0.06 3.465 0.535 3.405 0.535 3.405 0.06 3.055 0.06 3.055 0.535 2.995 0.535 2.995 0.06 2.645 0.06 2.645 0.535 2.585 0.535 2.585 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
  END VSS
  PIN ISOn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06435 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.911422 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.355 0.67 3.645 0.79 ;
    END
  END ISOn
  OBS
    LAYER Metal1 ;
      POLYGON 3.705 2.66 3.24 2.66 3.24 3.04 3.18 3.04 3.18 2.66 2.83 2.66 2.83 3.04 2.77 3.04 2.77 2.45 2.2 2.45 2.2 1.99 2.26 1.99 2.26 2.39 2.71 2.39 2.71 2.37 2.83 2.37 2.83 2.6 3.705 2.6 ;
      POLYGON 3.635 3.245 0.84 3.245 0.84 2.95 0.9 2.95 0.9 3.185 1.69 3.185 1.69 1.925 1.75 1.925 1.75 3.185 2.155 3.185 2.155 2.78 2.215 2.78 2.215 3.185 2.565 3.185 2.565 2.78 2.625 2.78 2.625 3.185 2.975 3.185 2.975 2.78 3.035 2.78 3.035 3.185 3.575 3.185 3.575 2.78 3.635 2.78 ;
      POLYGON 3.53 1.57 3.405 1.57 3.405 0.96 3.465 0.96 3.465 1.51 3.53 1.51 ;
      POLYGON 3.26 0.705 1.75 0.705 1.75 1.465 1.69 1.465 1.69 0.645 2.79 0.645 2.79 0.275 2.85 0.275 2.85 0.645 3.2 0.645 3.2 0.275 3.26 0.275 ;
      POLYGON 2.73 2.21 2.415 2.21 2.415 2.15 2.67 2.15 2.67 1.99 2.73 1.99 ;
      POLYGON 2.42 3.04 2.36 3.04 2.36 2.66 2.01 2.66 2.01 3.04 1.95 3.04 1.95 2.275 2.01 2.275 2.01 2.6 2.42 2.6 ;
      POLYGON 1.575 2.74 1.515 2.74 1.515 3.01 1.105 3.01 1.105 3.095 1.045 3.095 1.045 2.95 1.455 2.95 1.455 2.19 1.045 2.19 1.045 1.975 1.105 1.975 1.105 2.13 1.515 2.13 1.515 2.68 1.575 2.68 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSLH_ISONH_X1_TO_ON

MACRO LSLH_ISONL_X1_FROM_OFF
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSLH_ISONL_X1_FROM_OFF 0 0 ;
  SIZE 4 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 0.295 1.77 0.295 2.255 0.235 2.255 0.235 1.77 0 1.77 0 1.65 4 1.65 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0513 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.22 2.68 0.365 2.82 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.881875 LAYER Metal1 ;
    ANTENNADIFFAREA 2.0298 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0837 LAYER Metal1 ;
      ANTENNAMAXAREACAR 34.4310035 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 257.0250895 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.38 2.465 3.235 2.465 3.235 3.185 3.175 3.185 3.175 1.955 3.235 1.955 3.235 2.09 3.38 2.09 ;
    END
  END Y
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.03 2.345 2.97 2.345 2.97 2.265 2.645 2.265 2.645 2.49 2.765 2.49 2.765 2.63 2.435 2.63 2.435 2.49 2.585 2.49 2.585 2.265 2.27 2.265 2.27 1.93 1.45 1.93 1.45 2.265 1.39 2.265 1.39 1.87 2.33 1.87 2.33 2.205 2.585 2.205 2.585 2 2.645 2 2.645 2.205 2.97 2.205 2.97 1.955 3.03 1.955 ;
    END
  END ExtVDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 3.48 0 3.48 0 3.36 2.97 3.36 2.97 2.925 3.03 2.925 3.03 3.36 4 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.015 0.06 3.015 0.51 2.955 0.51 2.955 0.06 2.605 0.06 2.605 0.51 2.545 0.51 2.545 0.06 2.195 0.06 2.195 0.51 2.135 0.51 2.135 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
  END VSS
  PIN ISOn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.068175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.8261825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.68 0.79 2.965 0.92 ;
    END
  END ISOn
  OBS
    LAYER Metal1 ;
      POLYGON 3.165 1.545 2.79 1.545 2.79 1.045 2.85 1.045 2.85 1.485 3.165 1.485 ;
      POLYGON 3.09 2.76 3.06 2.76 3.06 2.79 2.635 2.79 2.635 3.13 2.575 3.13 2.575 2.79 2.225 2.79 2.225 3.13 2.165 3.13 2.165 2.53 1.595 2.53 1.595 2.05 1.655 2.05 1.655 2.47 2.265 2.47 2.265 2.53 2.225 2.53 2.225 2.73 2.97 2.73 2.97 2.7 3.09 2.7 ;
      POLYGON 2.81 0.72 0.99 0.72 0.99 1.515 0.93 1.515 0.93 0.66 2.34 0.66 2.34 0.25 2.4 0.25 2.4 0.66 2.75 0.66 2.75 0.25 2.81 0.25 ;
      RECT 2.585 1.045 2.645 1.575 ;
      POLYGON 2.43 3.255 0.235 3.255 0.235 2.98 0.295 2.98 0.295 3.195 0.93 3.195 0.93 1.97 0.99 1.97 0.99 3.195 1.55 3.195 1.55 2.87 1.61 2.87 1.61 3.195 1.96 3.195 1.96 2.87 2.02 2.87 2.02 3.195 2.37 3.195 2.37 2.87 2.43 2.87 ;
      POLYGON 2.125 2.39 1.81 2.39 1.81 2.33 2.065 2.33 2.065 2.05 2.125 2.05 ;
      POLYGON 1.815 3.13 1.755 3.13 1.755 2.74 1.405 2.74 1.405 3.13 1.345 3.13 1.345 2.335 1.405 2.335 1.405 2.68 1.815 2.68 ;
      POLYGON 0.62 2.855 0.5 2.855 0.5 3.125 0.44 3.125 0.44 2.04 0.5 2.04 0.5 2.795 0.62 2.795 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSLH_ISONL_X1_FROM_OFF

MACRO LSLH_ISONL_X1_TO_ON
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSLH_ISONL_X1_TO_ON 0 0 ;
  SIZE 4 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 3.485 1.77 3.485 2.345 3.425 2.345 3.425 1.77 2.92 1.77 2.92 2.205 2.86 2.205 2.86 1.77 2.04 1.77 2.04 2.205 1.98 2.205 1.98 1.77 0 1.77 0 1.65 3.185 1.65 3.185 1.185 3.245 1.185 3.245 1.65 4 1.65 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0513 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.16374275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.61 2.69 0.84 2.83 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.78745 LAYER Metal1 ;
    ANTENNADIFFAREA 2.0298 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0837 LAYER Metal1 ;
      ANTENNAMAXAREACAR 33.3028675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 247.09677425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.78 2.635 3.69 2.635 3.69 3.185 3.63 3.185 3.63 1.955 3.69 1.955 3.69 2.29 3.78 2.29 ;
    END
  END Y
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.165 2.63 0.775 2.63 0.775 2.49 0.825 2.49 0.825 1.975 0.885 1.975 0.885 2.49 1.165 2.49 ;
    END
  END ExtVDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 3.48 0 3.48 0 3.36 3.425 3.36 3.425 2.925 3.485 2.925 3.485 3.36 4 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.45 0.06 3.45 0.535 3.39 0.535 3.39 0.06 3.04 0.06 3.04 0.535 2.98 0.535 2.98 0.06 2.63 0.06 2.63 0.535 2.57 0.535 2.57 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
  END VSS
  PIN ISOn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.056475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.124834 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.295 0.975 3.565 1.105 ;
    END
  END ISOn
  OBS
    LAYER Metal1 ;
      POLYGON 3.56 2.53 3.225 2.53 3.225 3.04 3.165 3.04 3.165 2.53 2.815 2.53 2.815 3.04 2.755 3.04 2.755 2.45 2.185 2.45 2.185 1.99 2.245 1.99 2.245 2.39 2.695 2.39 2.695 2.37 2.815 2.37 2.815 2.47 3.56 2.47 ;
      POLYGON 3.55 1.585 3.49 1.585 3.49 1.505 3.39 1.505 3.39 1.185 3.45 1.185 3.45 1.445 3.55 1.445 ;
      POLYGON 3.245 0.8 1.735 0.8 1.735 1.465 1.675 1.465 1.675 0.74 2.775 0.74 2.775 0.275 2.835 0.275 2.835 0.74 3.185 0.74 3.185 0.275 3.245 0.275 ;
      POLYGON 3.02 3.245 0.825 3.245 0.825 2.95 0.885 2.95 0.885 3.185 1.675 3.185 1.675 1.925 1.735 1.925 1.735 3.185 2.14 3.185 2.14 2.78 2.2 2.78 2.2 3.185 2.55 3.185 2.55 2.78 2.61 2.78 2.61 3.185 2.96 3.185 2.96 2.78 3.02 2.78 ;
      POLYGON 2.715 2.21 2.4 2.21 2.4 2.15 2.655 2.15 2.655 1.99 2.715 1.99 ;
      POLYGON 2.405 3.04 2.345 3.04 2.345 2.66 1.995 2.66 1.995 3.04 1.935 3.04 1.935 2.275 1.995 2.275 1.995 2.6 2.405 2.6 ;
      POLYGON 1.56 2.74 1.5 2.74 1.5 3.01 1.09 3.01 1.09 3.095 1.03 3.095 1.03 2.95 1.44 2.95 1.44 2.19 1.03 2.19 1.03 1.975 1.09 1.975 1.09 2.13 1.5 2.13 1.5 2.68 1.56 2.68 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSLH_ISONL_X1_TO_ON

MACRO LSLHX1_FROM
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSLHX1_FROM 0 0 ;
  SIZE 4 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 0.295 1.77 0.295 2.255 0.235 2.255 0.235 1.77 0 1.77 0 1.65 4 1.65 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0513 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.6959065 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.22 2.675 0.365 2.82 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.80635 LAYER Metal1 ;
    ANTENNADIFFAREA 1.292 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0837 LAYER Metal1 ;
      ANTENNAMAXAREACAR 21.5812425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 158.27957 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.19 3.185 3.13 3.185 3.13 2.51 3.02 2.51 3.02 2.305 3.065 2.305 3.065 1.955 3.125 1.955 3.125 2.305 3.19 2.305 ;
    END
  END Y
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.92 2.345 2.86 2.345 2.86 2.265 2.645 2.265 2.645 2.49 2.765 2.49 2.765 2.63 2.435 2.63 2.435 2.49 2.585 2.49 2.585 2.265 2.27 2.265 2.27 1.93 1.45 1.93 1.45 2.265 1.39 2.265 1.39 1.87 2.33 1.87 2.33 2.205 2.86 2.205 2.86 1.955 2.92 1.955 ;
    END
  END ExtVDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 3.48 0 3.48 0 3.36 0.235 3.36 0.235 2.98 0.295 2.98 0.295 3.36 1.55 3.36 1.55 2.925 1.61 2.925 1.61 3.36 1.96 3.36 1.96 2.925 2.02 2.925 2.02 3.36 2.37 3.36 2.37 2.925 2.43 2.925 2.43 3.36 2.97 3.36 2.97 3.185 2.925 3.185 2.925 2.925 2.985 2.925 2.985 3.125 3.03 3.125 3.03 3.36 4 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 4 0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.045 2.815 2.635 2.815 2.635 3.185 2.575 3.185 2.575 2.815 2.225 2.815 2.225 3.185 2.165 3.185 2.165 2.53 1.595 2.53 1.595 2.05 1.655 2.05 1.655 2.47 2.225 2.47 2.225 2.755 3.045 2.755 ;
      POLYGON 2.125 2.39 1.81 2.39 1.81 2.33 2.065 2.33 2.065 2.05 2.125 2.05 ;
      POLYGON 1.815 3.185 1.755 3.185 1.755 2.815 1.405 2.815 1.405 3.185 1.345 3.185 1.345 2.335 1.405 2.335 1.405 2.755 1.815 2.755 ;
      POLYGON 0.62 2.885 0.5 2.885 0.5 3.125 0.44 3.125 0.44 2.04 0.5 2.04 0.5 2.825 0.62 2.825 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSLHX1_FROM

MACRO LSLHX1_TO
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LSLHX1_TO 0 0 ;
  SIZE 4 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 3.63 1.77 3.63 2.345 3.57 2.345 3.57 1.77 2.93 1.77 2.93 2.265 2.87 2.265 2.87 1.77 2.05 1.77 2.05 2.265 1.99 2.265 1.99 1.77 0 1.77 0 1.65 4 1.65 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0513 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.27485375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.93 2.9 0.875 2.9 0.875 3.01 0.6 3.01 0.6 2.78 0.93 2.78 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.827825 LAYER Metal1 ;
    ANTENNADIFFAREA 1.3512 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0837 LAYER Metal1 ;
      ANTENNAMAXAREACAR 21.8378135 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 159.24731175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.94 2.635 3.835 2.635 3.835 3.185 3.775 3.185 3.775 1.955 3.835 1.955 3.835 2.49 3.94 2.49 ;
    END
  END Y
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 2.63 0.815 2.63 0.815 2.49 0.945 2.49 0.945 1.975 1.005 1.975 1.005 2.49 1.4 2.49 ;
    END
  END ExtVDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 3.48 0 3.48 0 3.36 0.945 3.36 0.945 3.03 1.005 3.03 1.005 3.36 2.15 3.36 2.15 2.925 2.21 2.925 2.21 3.36 2.56 3.36 2.56 2.925 2.62 2.925 2.62 3.36 2.97 3.36 2.97 2.925 3.03 2.925 3.03 3.36 3.57 3.36 3.57 2.925 3.63 2.925 3.63 3.36 4 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 4 0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.69 2.785 3.235 2.785 3.235 3.185 3.175 3.185 3.175 2.785 2.825 2.785 2.825 3.185 2.765 3.185 2.765 2.53 2.195 2.53 2.195 2.05 2.255 2.05 2.255 2.47 2.825 2.47 2.825 2.725 3.69 2.725 ;
      POLYGON 2.725 2.39 2.41 2.39 2.41 2.33 2.665 2.33 2.665 2.05 2.725 2.05 ;
      POLYGON 2.415 3.185 2.355 3.185 2.355 2.815 2.005 2.815 2.005 3.185 1.945 3.185 1.945 2.335 2.005 2.335 2.005 2.755 2.415 2.755 ;
      POLYGON 1.775 2.885 1.715 2.885 1.715 3.09 1.21 3.09 1.21 3.175 1.15 3.175 1.15 3.03 1.655 3.03 1.655 2.19 1.15 2.19 1.15 1.975 1.21 1.975 1.21 2.13 1.715 2.13 1.715 2.825 1.775 2.825 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END LSLHX1_TO

MACRO MDFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MDFFHQX1 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.616225 LAYER Metal1 ;
    ANTENNADIFFAREA 3.24895 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2601 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.05853525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 79.25605525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.2 1.475 0.14 1.475 0.14 0.73 0.06 0.73 0.06 0.6 0.14 0.6 0.14 0.54 0.2 0.54 ;
    END
  END Q
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.88778875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.77 0.745 4.71 0.745 4.71 0.705 3.995 0.705 3.995 0.945 3.935 0.945 3.935 0.645 4.635 0.645 4.635 0.625 4.77 0.625 ;
    END
  END S0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.61 0.895 4.565 0.895 4.565 1.04 4.265 1.04 4.265 0.805 4.61 0.805 ;
    END
  END D1
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.675 0.91 3.595 0.91 3.595 0.73 3.46 0.73 3.46 0.545 3.54 0.545 3.54 0.65 3.675 0.65 ;
    END
  END D0
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.565 1.035 0.54 1.035 0.54 1.255 0.46 1.255 0.46 0.79 0.485 0.79 0.485 0.78 0.565 0.78 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 1.77 0 1.77 0 1.65 0.345 1.65 0.345 1.355 0.405 1.355 0.405 1.65 1.11 1.65 1.11 1.29 1.23 1.29 1.23 1.35 1.17 1.35 1.17 1.65 2.365 1.65 2.365 1.365 2.485 1.365 2.485 1.425 2.425 1.425 2.425 1.65 3.615 1.65 3.615 1.17 3.675 1.17 3.675 1.65 4.425 1.65 4.425 1.315 4.485 1.315 4.485 1.65 5 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 0.06 4.54 0.06 4.54 0.525 4.48 0.525 4.48 0.06 3.675 0.06 3.675 0.415 3.615 0.415 3.615 0.06 2.425 0.06 2.425 0.19 2.485 0.19 2.485 0.25 2.365 0.25 2.365 0.06 1.225 0.06 1.225 0.49 1.165 0.49 1.165 0.06 0.405 0.06 0.405 0.52 0.345 0.52 0.345 0.06 0 0.06 0 -0.06 5 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.93 1.2 4.845 1.2 4.845 1.26 4.785 1.26 4.785 1.2 4.105 1.2 4.105 0.885 4.165 0.885 4.165 1.14 4.87 1.14 4.87 0.43 4.93 0.43 ;
      POLYGON 4.23 0.545 3.835 0.545 3.835 1.045 4.005 1.045 4.005 1.435 3.945 1.435 3.945 1.105 3.775 1.105 3.775 1.07 3.21 1.07 3.21 1.13 3.15 1.13 3.15 1.01 3.21 1.01 3.21 0.545 3.15 0.545 3.15 0.485 3.27 0.485 3.27 1.01 3.775 1.01 3.775 0.485 4.17 0.485 4.17 0.425 4.23 0.425 ;
      POLYGON 3.47 1.23 3.37 1.23 3.37 1.29 2.99 1.29 2.99 0.355 2.67 0.355 2.67 0.615 2.73 0.615 2.73 0.735 2.67 0.735 2.67 0.675 2.61 0.675 2.61 0.41 2.205 0.41 2.205 0.385 1.885 0.385 1.885 0.66 1.87 0.66 1.87 0.81 1.585 0.81 1.585 0.87 1.525 0.87 1.525 0.75 1.81 0.75 1.81 0.615 1.825 0.615 1.825 0.325 2.265 0.325 2.265 0.35 2.61 0.35 2.61 0.295 3.44 0.295 3.44 0.415 3.38 0.415 3.38 0.355 3.05 0.355 3.05 1.23 3.31 1.23 3.31 1.17 3.47 1.17 ;
      POLYGON 2.89 1.205 2.83 1.205 2.83 1.005 2.29 1.005 2.29 0.755 2.35 0.755 2.35 0.945 2.83 0.945 2.83 0.515 2.77 0.515 2.77 0.455 2.89 0.455 ;
      POLYGON 2.78 1.365 2.66 1.365 2.66 1.265 1.43 1.265 1.43 1.19 0.725 1.19 0.725 1.38 0.665 1.38 0.665 0.54 0.725 0.54 0.725 1.13 1.49 1.13 1.49 1.205 1.97 1.205 1.97 0.765 2.03 0.765 2.03 1.205 2.72 1.205 2.72 1.305 2.78 1.305 ;
      POLYGON 2.51 0.845 2.45 0.845 2.45 0.655 2.19 0.655 2.19 1.105 2.13 1.105 2.13 0.57 1.985 0.57 1.985 0.485 2.105 0.485 2.105 0.51 2.19 0.51 2.19 0.595 2.51 0.595 ;
      POLYGON 1.725 0.545 1.425 0.545 1.425 0.97 1.65 0.97 1.65 1.105 1.59 1.105 1.59 1.03 1.045 1.03 1.045 0.87 1.035 0.87 1.035 0.75 1.105 0.75 1.105 0.97 1.365 0.97 1.365 0.485 1.725 0.485 ;
      POLYGON 1.265 0.865 1.205 0.865 1.205 0.65 0.885 0.65 0.885 0.97 0.945 0.97 0.945 1.03 0.825 1.03 0.825 0.44 0.565 0.44 0.565 0.68 0.36 0.68 0.36 0.82 0.3 0.82 0.3 0.62 0.505 0.62 0.505 0.38 1.02 0.38 1.02 0.59 1.265 0.59 ;
  END
END MDFFHQX1

MACRO MDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MDFFHQX2 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.763325 LAYER Metal1 ;
    ANTENNADIFFAREA 3.4928 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.28935 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.55011225 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 74.88335925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.36 1.335 0.3 1.335 0.3 0.92 0.26 0.92 0.26 0.79 0.3 0.79 0.3 0.54 0.36 0.54 ;
    END
  END Q
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 12.2442245 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.165 0.895 5.035 0.895 5.035 0.875 5.025 0.875 5.025 0.815 5.085 0.815 5.085 0.56 4.56 0.56 4.56 0.67 4.44 0.67 4.44 0.56 4.255 0.56 4.255 0.88 4.195 0.88 4.195 0.5 5.145 0.5 5.145 0.815 5.165 0.815 ;
    END
  END S0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.925 0.975 4.66 0.975 4.66 0.785 4.845 0.785 4.845 0.66 4.925 0.66 ;
    END
  END D1
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.935 0.805 3.855 0.805 3.855 0.73 3.66 0.73 3.66 0.5 3.74 0.5 3.74 0.645 3.935 0.645 ;
    END
  END D0
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.815 1.02 0.54 1.02 0.54 1.115 0.46 1.115 0.46 0.94 0.635 0.94 0.635 0.89 0.815 0.89 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 1.77 0 1.77 0 1.65 0.095 1.65 0.095 1.02 0.155 1.02 0.155 1.65 0.505 1.65 0.505 1.215 0.565 1.215 0.565 1.65 1.34 1.65 1.34 1.28 1.4 1.28 1.4 1.65 2.615 1.65 2.615 1.28 2.735 1.28 2.735 1.34 2.675 1.34 2.675 1.65 3.875 1.65 3.875 1.065 3.935 1.065 3.935 1.65 4.675 1.65 4.675 1.25 4.735 1.25 4.735 1.65 5.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 0.06 4.795 0.06 4.795 0.4 4.735 0.4 4.735 0.06 3.935 0.06 3.935 0.4 3.875 0.4 3.875 0.06 2.735 0.06 2.735 0.25 2.615 0.25 2.615 0.19 2.675 0.19 2.675 0.06 1.425 0.06 1.425 0.445 1.365 0.445 1.365 0.06 0.565 0.06 0.565 0.52 0.505 0.52 0.505 0.06 0.155 0.06 0.155 0.52 0.095 0.52 0.095 0.06 0 0.06 0 -0.06 5.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.325 1.135 5.19 1.135 5.19 1.195 5.13 1.195 5.13 1.135 4.43 1.135 4.43 0.82 4.49 0.82 4.49 1.075 5.265 1.075 5.265 0.715 5.245 0.715 5.245 0.42 5.305 0.42 5.305 0.655 5.325 0.655 ;
      POLYGON 4.48 0.4 4.095 0.4 4.095 0.98 4.33 0.98 4.33 1.37 4.27 1.37 4.27 1.04 4.035 1.04 4.035 0.965 3.5 0.965 3.5 1.04 3.44 1.04 3.44 0.44 3.56 0.44 3.56 0.5 3.5 0.5 3.5 0.905 4.035 0.905 4.035 0.34 4.42 0.34 4.42 0.28 4.48 0.28 ;
      POLYGON 3.73 0.4 3.67 0.4 3.67 0.34 3.34 0.34 3.34 1.185 3.73 1.185 3.73 1.245 3.28 1.245 3.28 0.34 2.96 0.34 2.96 0.6 3.02 0.6 3.02 0.66 2.9 0.66 2.9 0.41 2.455 0.41 2.455 0.34 2.135 0.34 2.135 0.645 2.07 0.645 2.07 0.765 1.785 0.765 1.785 0.825 1.725 0.825 1.725 0.705 2.01 0.705 2.01 0.585 2.075 0.585 2.075 0.28 2.515 0.28 2.515 0.35 2.9 0.35 2.9 0.28 3.73 0.28 ;
      POLYGON 3.18 1.18 3.12 1.18 3.12 0.82 2.51 0.82 2.51 0.76 3.12 0.76 3.12 0.5 3.06 0.5 3.06 0.44 3.18 0.44 ;
      POLYGON 3.07 1.34 2.95 1.34 2.95 1.18 2.25 1.18 2.25 1.205 1.63 1.205 1.63 1.18 0.77 1.18 0.77 1.24 0.71 1.24 0.71 1.12 0.915 1.12 0.915 0.54 0.975 0.54 0.975 1.12 1.69 1.12 1.69 1.145 2.19 1.145 2.19 0.74 2.25 0.74 2.25 1.12 3.01 1.12 3.01 1.28 3.07 1.28 ;
      POLYGON 2.8 0.66 2.41 0.66 2.41 1.02 2.35 1.02 2.35 0.57 2.235 0.57 2.235 0.44 2.355 0.44 2.355 0.51 2.41 0.51 2.41 0.6 2.8 0.6 ;
      POLYGON 1.975 0.485 1.91 0.485 1.91 0.605 1.625 0.605 1.625 0.925 1.85 0.925 1.85 1.045 1.79 1.045 1.79 0.985 1.245 0.985 1.245 0.84 1.235 0.84 1.235 0.72 1.305 0.72 1.305 0.925 1.565 0.925 1.565 0.545 1.85 0.545 1.85 0.425 1.975 0.425 ;
      POLYGON 1.465 0.82 1.405 0.82 1.405 0.605 1.135 0.605 1.135 0.9 1.145 0.9 1.145 1.02 1.085 1.02 1.085 0.94 1.075 0.94 1.075 0.44 0.815 0.44 0.815 0.79 0.46 0.79 0.46 0.73 0.755 0.73 0.755 0.38 1.22 0.38 1.22 0.545 1.465 0.545 ;
  END
END MDFFHQX2

MACRO MDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MDFFHQX4 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.60066 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.165 0.715 4.53 0.715 4.53 0.93 4.47 0.93 4.47 0.655 5.035 0.655 5.035 0.625 5.165 0.625 ;
    END
  END S0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.20512825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.82 0.815 5.06 0.985 ;
    END
  END D1
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.21 0.93 4.13 0.93 4.13 0.92 3.86 0.92 3.86 0.79 3.94 0.79 3.94 0.84 4.13 0.84 4.13 0.75 4.21 0.75 ;
    END
  END D0
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.69 0.34 1.19 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8383 LAYER Metal1 ;
    ANTENNADIFFAREA 3.66465 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.371025 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.64988875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 60.0283 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.065 1.075 0.46 1.075 0.46 0.79 0.525 0.79 0.525 0.54 0.585 0.54 0.585 0.85 0.54 0.85 0.54 1.015 1.005 1.015 1.005 0.54 1.065 0.54 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 1.77 0 1.77 0 1.65 0.27 1.65 0.27 1.51 0.33 1.51 0.33 1.65 0.71 1.65 0.71 1.45 0.83 1.45 0.83 1.51 0.77 1.51 0.77 1.65 1.18 1.65 1.18 1.45 1.3 1.45 1.3 1.51 1.24 1.51 1.24 1.65 1.65 1.65 1.65 1.45 1.77 1.45 1.77 1.51 1.71 1.51 1.71 1.65 2.85 1.65 2.85 1.4 2.97 1.4 2.97 1.46 2.91 1.46 2.91 1.65 4.19 1.65 4.19 1.26 4.25 1.26 4.25 1.65 4.915 1.65 4.915 1.26 4.975 1.26 4.975 1.65 5.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 0.06 5.05 0.06 5.05 0.525 4.99 0.525 4.99 0.06 4.18 0.06 4.18 0.55 4.12 0.55 4.12 0.06 2.97 0.06 2.97 0.255 2.85 0.255 2.85 0.195 2.91 0.195 2.91 0.06 1.71 0.06 1.71 0.52 1.65 0.52 1.65 0.06 1.29 0.06 1.29 0.52 1.23 0.52 1.23 0.06 0.79 0.06 0.79 0.52 0.73 0.52 0.73 0.06 0.38 0.06 0.38 0.52 0.32 0.52 0.32 0.06 0 0.06 0 -0.06 5.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.325 1.145 5.255 1.145 5.255 1.205 5.195 1.205 5.195 1.145 4.66 1.145 4.66 0.83 4.72 0.83 4.72 1.085 5.265 1.085 5.265 0.43 5.325 0.43 ;
      POLYGON 4.74 0.555 4.37 0.555 4.37 1.03 4.56 1.03 4.56 1.38 4.5 1.38 4.5 1.09 3.625 1.09 3.625 1.03 3.685 1.03 3.685 0.515 3.805 0.515 3.805 0.575 3.745 0.575 3.745 1.03 4.31 1.03 4.31 0.495 4.68 0.495 4.68 0.435 4.74 0.435 ;
      POLYGON 4.075 1.255 3.465 1.255 3.465 0.81 3.525 0.81 3.525 0.415 3.205 0.415 3.205 0.775 3.145 0.775 3.145 0.415 2.37 0.415 2.37 0.725 2.335 0.725 2.335 0.785 2.07 0.785 2.07 0.905 2.01 0.905 2.01 0.725 2.275 0.725 2.275 0.665 2.31 0.665 2.31 0.355 3.975 0.355 3.975 0.55 3.915 0.55 3.915 0.415 3.585 0.415 3.585 0.93 3.525 0.93 3.525 1.195 4.075 1.195 ;
      POLYGON 3.425 0.575 3.365 0.575 3.365 1.265 3.305 1.265 3.305 0.935 2.765 0.935 2.765 0.845 2.885 0.845 2.885 0.875 3.305 0.875 3.305 0.515 3.425 0.515 ;
      POLYGON 3.255 1.425 3.135 1.425 3.135 1.3 2.505 1.3 2.505 1.35 0.085 1.35 0.085 0.54 0.145 0.54 0.145 1.29 2.445 1.29 2.445 0.8 2.505 0.8 2.505 1.24 3.195 1.24 3.195 1.365 3.255 1.365 ;
      POLYGON 3.045 0.745 2.665 0.745 2.665 1.14 2.605 1.14 2.605 0.575 2.47 0.575 2.47 0.515 2.665 0.515 2.665 0.685 3.045 0.685 ;
      POLYGON 2.21 0.565 1.91 0.565 1.91 1.005 2.145 1.005 2.145 1.19 2.085 1.19 2.085 1.065 1.85 1.065 1.85 0.925 1.52 0.925 1.52 0.805 1.58 0.805 1.58 0.865 1.85 0.865 1.85 0.505 2.21 0.505 ;
      POLYGON 1.75 0.765 1.69 0.765 1.69 0.705 1.42 0.705 1.42 1.025 1.535 1.025 1.535 1.085 1.36 1.085 1.36 0.705 1.225 0.705 1.225 0.82 1.165 0.82 1.165 0.645 1.445 0.645 1.445 0.485 1.505 0.485 1.505 0.645 1.75 0.645 ;
  END
END MDFFHQX4

MACRO MDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MDFFHQX8 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.21782175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 0.745 6.34 0.745 6.34 0.705 5.685 0.705 5.685 0.755 5.595 0.755 5.595 0.965 5.535 0.965 5.535 0.695 5.625 0.695 5.625 0.645 6.235 0.645 6.235 0.625 6.4 0.625 ;
    END
  END S0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.24 0.885 6.165 0.885 6.165 1.01 5.865 1.01 5.865 0.805 6.24 0.805 ;
    END
  END D1
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.275 1.015 5.195 1.015 5.195 0.92 5.06 0.92 5.06 0.65 5.14 0.65 5.14 0.79 5.275 0.79 ;
    END
  END D0
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.83 0.895 2.555 0.895 2.555 0.815 2.72 0.815 2.72 0.59 2.83 0.59 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6952 LAYER Metal1 ;
    ANTENNADIFFAREA 4.57105 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.528525 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.991533 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 54.8034625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.36 0.65 1.315 0.65 1.315 0.9 1.36 0.9 1.36 1.345 1.3 1.345 1.3 0.96 1.255 0.96 1.255 0.8 0.95 0.8 0.95 1.345 0.89 1.345 0.89 0.73 0.54 0.73 0.54 1.345 0.48 1.345 0.48 0.73 0.13 0.73 0.13 1.345 0.07 1.345 0.07 0.73 0.06 0.73 0.06 0.6 0.07 0.6 0.07 0.54 0.14 0.54 0.14 0.67 0.48 0.67 0.48 0.54 0.54 0.54 0.54 0.67 0.89 0.67 0.89 0.54 0.95 0.54 0.95 0.74 1.255 0.74 1.255 0.59 1.3 0.59 1.3 0.53 1.36 0.53 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 1.77 0 1.77 0 1.65 0.275 1.65 0.275 0.9 0.335 0.9 0.335 1.65 0.685 1.65 0.685 0.9 0.745 0.9 0.745 1.65 1.095 1.65 1.095 0.9 1.155 0.9 1.155 1.65 1.505 1.65 1.505 0.905 1.565 0.905 1.565 1.65 1.945 1.65 1.945 1.055 2.005 1.055 2.005 1.65 2.93 1.65 2.93 1.51 2.99 1.51 2.99 1.65 4.055 1.65 4.055 1.315 4.175 1.315 4.175 1.375 4.115 1.375 4.115 1.65 5.235 1.65 5.235 1.285 5.295 1.285 5.295 1.65 6.055 1.65 6.055 1.285 6.115 1.285 6.115 1.65 6.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 0.06 6.115 0.06 6.115 0.525 6.055 0.525 6.055 0.06 5.365 0.06 5.365 0.435 5.305 0.435 5.305 0.06 4.175 0.06 4.175 0.17 4.055 0.17 4.055 0.06 2.915 0.06 2.915 0.17 2.795 0.17 2.795 0.06 1.975 0.06 1.975 0.485 1.915 0.485 1.915 0.06 1.565 0.06 1.565 0.485 1.505 0.485 1.505 0.06 1.155 0.06 1.155 0.485 1.095 0.485 1.095 0.06 0.745 0.06 0.745 0.485 0.685 0.485 0.685 0.06 0.335 0.06 0.335 0.485 0.275 0.485 0.275 0.06 0 0.06 0 -0.06 6.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.56 1.17 6.35 1.17 6.35 1.23 6.29 1.23 6.29 1.17 5.705 1.17 5.705 0.855 5.765 0.855 5.765 1.11 6.5 1.11 6.5 0.525 6.29 0.525 6.29 0.405 6.35 0.405 6.35 0.465 6.56 0.465 ;
      POLYGON 5.805 0.545 5.525 0.545 5.525 0.595 5.435 0.595 5.435 1.115 5.605 1.115 5.605 1.405 5.545 1.405 5.545 1.175 4.84 1.175 4.84 0.98 4.9 0.98 4.9 0.515 4.84 0.515 4.84 0.455 4.96 0.455 4.96 1.115 5.375 1.115 5.375 0.535 5.465 0.535 5.465 0.485 5.745 0.485 5.745 0.425 5.805 0.425 ;
      POLYGON 5.13 0.55 5.07 0.55 5.07 0.355 4.74 0.355 4.74 1.315 5.12 1.315 5.12 1.375 4.68 1.375 4.68 0.355 4.36 0.355 4.36 0.615 4.41 0.615 4.41 0.735 4.3 0.735 4.3 0.355 3.575 0.355 3.575 0.615 3.69 0.615 3.69 0.735 3.63 0.735 3.63 0.675 3.515 0.675 3.515 0.295 5.13 0.295 ;
      POLYGON 4.58 1.215 4.52 1.215 4.52 0.895 4.01 0.895 4.01 0.855 3.95 0.855 3.95 0.795 4.07 0.795 4.07 0.835 4.52 0.835 4.52 0.515 4.46 0.515 4.46 0.455 4.58 0.455 ;
      POLYGON 4.47 1.375 4.35 1.375 4.35 1.215 3.09 1.215 3.09 0.49 2.455 0.49 2.455 0.995 2.705 0.995 2.705 1.115 2.645 1.115 2.645 1.055 2.395 1.055 2.395 0.43 3.15 0.43 3.15 1.155 3.47 1.155 3.47 0.835 3.41 0.835 3.41 0.775 3.53 0.775 3.53 1.155 4.41 1.155 4.41 1.315 4.47 1.315 ;
      POLYGON 4.2 0.715 4.14 0.715 4.14 0.695 3.85 0.695 3.85 1.055 3.79 1.055 3.79 0.515 3.675 0.515 3.675 0.455 3.85 0.455 3.85 0.635 4.14 0.635 4.14 0.595 4.2 0.595 ;
      POLYGON 3.37 1.055 3.31 1.055 3.31 0.995 3.25 0.995 3.25 0.33 2.135 0.33 2.135 0.795 2.075 0.795 2.075 0.27 3.31 0.27 3.31 0.935 3.37 0.935 ;
      POLYGON 2.99 1.275 2.21 1.275 2.21 1.345 2.15 1.345 2.15 0.955 1.8 0.955 1.8 1.345 1.74 1.345 1.74 0.955 1.71 0.955 1.71 0.805 1.415 0.805 1.415 0.745 1.71 0.745 1.71 0.505 1.77 0.505 1.77 0.895 2.235 0.895 2.235 0.505 2.295 0.505 2.295 1.215 2.93 1.215 2.93 0.74 2.99 0.74 ;
  END
END MDFFHQX8

MACRO MX2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8004 LAYER Metal1 ;
    ANTENNADIFFAREA 0.7575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXAREACAR 17.610561 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 134.85148525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.57 1.33 0.57 1.33 1.075 1.19 1.075 1.19 1.415 1.13 1.415 1.13 1.01 1.27 1.01 1.27 0.57 1.13 0.57 1.13 0.23 1.19 0.23 1.19 0.37 1.34 0.37 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.888889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.165 0.92 0.885 0.92 0.885 0.72 0.98 0.72 0.98 0.78 1.165 0.78 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.74 0.41 0.92 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.287037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.58 1.195 0.2 1.195 0.2 0.98 0.26 0.98 0.26 1.135 0.43 1.135 0.43 0.98 0.52 0.98 0.52 0.835 0.58 0.835 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.295 0.335 1.295 0.335 1.65 0.925 1.65 0.925 1.2 0.985 1.2 0.985 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 0.955 0.06 0.955 0.35 0.895 0.35 0.895 0.06 0.335 0.06 0.335 0.35 0.275 0.35 0.275 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.03 0.62 0.825 0.62 0.825 1.355 0.555 1.355 0.555 1.295 0.765 1.295 0.765 0.35 0.585 0.35 0.585 0.23 0.645 0.23 0.645 0.29 0.825 0.29 0.825 0.56 1.03 0.56 ;
      POLYGON 0.7 1.125 0.64 1.125 0.64 0.71 0.525 0.71 0.525 0.51 0.115 0.51 0.115 1.295 0.13 1.295 0.13 1.415 0.07 1.415 0.07 1.355 0.055 1.355 0.055 0.29 0.07 0.29 0.07 0.23 0.13 0.23 0.13 0.35 0.115 0.35 0.115 0.45 0.7 0.45 ;
  END
END MX2X1

MACRO MX2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8535 LAYER Metal1 ;
    ANTENNADIFFAREA 1.0052 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0747 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.42570275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 91.88755025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 0.73 1.66 0.73 1.66 0.66 1.56 0.66 1.56 1.105 1.525 1.105 1.525 1.435 1.465 1.435 1.465 1.045 1.5 1.045 1.5 0.485 1.465 0.485 1.465 0.365 1.525 0.365 1.525 0.425 1.56 0.425 1.56 0.6 1.74 0.6 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.895 1.3 0.895 1.3 1.215 1.22 1.215 1.22 0.815 1.4 0.815 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.62 1.035 0.44 1.035 0.44 0.955 0.46 0.955 0.46 0.635 0.54 0.635 0.54 0.955 0.62 0.955 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.074074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.215 0.26 1.215 0.26 0.98 0.34 0.98 0.34 1.135 0.72 1.135 0.72 0.93 0.8 0.93 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.41 1.65 0.41 1.315 0.47 1.315 0.47 1.65 1.26 1.65 1.26 1.315 1.32 1.315 1.32 1.65 1.67 1.65 1.67 1.045 1.73 1.045 1.73 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.73 0.06 1.73 0.375 1.67 0.375 1.67 0.06 1.32 0.06 1.32 0.375 1.26 0.375 1.26 0.06 0.47 0.06 0.47 0.375 0.41 0.375 0.41 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.4 0.645 1.12 0.645 1.12 1.335 0.89 1.335 0.89 1.275 1.06 1.275 1.06 0.375 0.735 0.375 0.735 0.255 0.795 0.255 0.795 0.315 1.12 0.315 1.12 0.585 1.4 0.585 ;
      POLYGON 0.96 1.155 0.9 1.155 0.9 0.805 0.64 0.805 0.64 0.535 0.16 0.535 0.16 1.315 0.265 1.315 0.265 1.435 0.205 1.435 0.205 1.375 0.1 1.375 0.1 0.475 0.205 0.475 0.205 0.28 0.265 0.28 0.265 0.475 0.76 0.475 0.76 0.745 0.96 0.745 ;
  END
END MX2X2

MACRO MX2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X4 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1918 LAYER Metal1 ;
    ANTENNADIFFAREA 1.505125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.140175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.50222925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 64.05564475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.995 0.53 1.63 0.53 1.63 0.98 1.74 0.98 1.74 1.05 1.995 1.05 1.995 1.48 1.935 1.48 1.935 1.11 1.585 1.11 1.585 1.48 1.525 1.48 1.525 1.05 1.57 1.05 1.57 0.48 1.495 0.48 1.495 0.42 1.63 0.42 1.63 0.47 1.935 0.47 1.935 0.39 1.995 0.39 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.47 0.895 1.315 0.895 1.315 1.105 1.18 1.105 1.18 0.95 1.235 0.95 1.235 0.815 1.47 0.815 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.63 0.54 1.13 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.039375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.60952375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 0.97 0.7 0.97 0.7 1.29 0.26 1.29 0.26 0.98 0.34 0.98 0.34 1.23 0.64 1.23 0.64 0.91 0.76 0.91 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 1.77 0 1.77 0 1.65 0.395 1.65 0.395 1.39 0.515 1.39 0.515 1.65 1.24 1.65 1.24 1.205 1.3 1.205 1.3 1.65 1.73 1.65 1.73 1.21 1.79 1.21 1.79 1.65 2.14 1.65 2.14 1.09 2.2 1.09 2.2 1.65 2.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 0.06 2.2 0.06 2.2 0.37 2.14 0.37 2.14 0.06 1.79 0.06 1.79 0.37 1.73 0.37 1.73 0.06 1.27 0.06 1.27 0.28 1.33 0.28 1.33 0.34 1.21 0.34 1.21 0.06 0.5 0.06 0.5 0.37 0.44 0.37 0.44 0.06 0 0.06 0 -0.06 2.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.47 0.715 1.08 0.715 1.08 1.265 0.87 1.265 0.87 1.325 0.81 1.325 0.81 1.205 1.02 1.205 1.02 0.37 0.87 0.37 0.87 0.25 0.93 0.25 0.93 0.31 1.08 0.31 1.08 0.655 1.47 0.655 ;
      POLYGON 0.92 1.105 0.86 1.105 0.86 0.66 0.8 0.66 0.8 0.53 0.16 0.53 0.16 1.39 0.295 1.39 0.295 1.45 0.1 1.45 0.1 0.47 0.205 0.47 0.205 0.335 0.265 0.335 0.265 0.47 0.92 0.47 ;
  END
END MX2X4

MACRO MX2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X6 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3599 LAYER Metal1 ;
    ANTENNADIFFAREA 1.815075 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.198675 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.844847 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 53.7561345 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.515 1.395 2.455 1.395 2.455 0.985 2.41 0.985 2.41 0.66 2.105 0.66 2.105 1.395 2.045 1.395 2.045 0.66 1.74 0.66 1.74 0.88 1.695 0.88 1.695 1.395 1.635 1.395 1.635 0.83 1.655 0.83 1.655 0.415 1.61 0.415 1.61 0.295 1.67 0.295 1.67 0.355 1.715 0.355 1.715 0.6 2.02 0.6 2.02 0.235 2.08 0.235 2.08 0.6 2.41 0.6 2.41 0.485 2.43 0.485 2.43 0.235 2.49 0.235 2.49 0.545 2.47 0.545 2.47 0.925 2.515 0.925 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.675 1.34 1.175 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 0.995 0.46 0.995 0.46 0.79 0.58 0.79 0.58 0.615 0.66 0.615 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.039375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.7714285 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.84 1.175 0.28 1.175 0.28 1.11 0.26 1.11 0.26 0.915 0.36 0.915 0.36 1.095 0.76 1.095 0.76 0.915 0.84 0.915 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 1.77 0 1.77 0 1.65 0.375 1.65 0.375 1.275 0.435 1.275 0.435 1.65 1.43 1.65 1.43 1.275 1.49 1.275 1.49 1.65 1.84 1.65 1.84 0.925 1.9 0.925 1.9 1.65 2.25 1.65 2.25 0.925 2.31 0.925 2.31 1.65 2.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 0.06 2.285 0.06 2.285 0.5 2.225 0.5 2.225 0.06 1.875 0.06 1.875 0.5 1.815 0.5 1.815 0.06 1.395 0.06 1.395 0.355 1.335 0.355 1.335 0.06 0.585 0.06 0.585 0.355 0.525 0.355 0.525 0.06 0 0.06 0 -0.06 2.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.555 0.73 1.495 0.73 1.495 0.575 1.16 0.575 1.16 1.18 1 1.18 1 1.24 0.94 1.24 0.94 1.12 1.1 1.12 1.1 0.355 0.835 0.355 0.835 0.235 0.895 0.235 0.895 0.295 1.16 0.295 1.16 0.515 1.555 0.515 ;
      POLYGON 1 1.02 0.94 1.02 0.94 0.815 0.77 0.815 0.77 0.515 0.16 0.515 0.16 1.18 0.18 1.18 0.18 1.3 0.12 1.3 0.12 1.23 0.1 1.23 0.1 0.455 0.225 0.455 0.225 0.32 0.285 0.32 0.285 0.455 0.83 0.455 0.83 0.755 1 0.755 ;
  END
END MX2X6

MACRO MX2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2X8 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.645175 LAYER Metal1 ;
    ANTENNADIFFAREA 2.34975 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.256275 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.41956875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 49.11911025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.325 1.435 3.265 1.435 3.265 1.05 2.915 1.05 2.915 1.435 2.855 1.435 2.855 1.05 2.505 1.05 2.505 1.435 2.445 1.435 2.445 1.05 2.14 1.05 2.14 1.11 2.095 1.11 2.095 1.435 2.035 1.435 2.035 0.99 2.06 0.99 2.06 0.59 2 0.59 2 0.53 2.12 0.53 2.12 0.98 2.14 0.98 2.14 0.99 3.265 0.99 3.265 0.615 2.49 0.615 2.49 0.6 2.415 0.6 2.415 0.54 2.535 0.54 2.535 0.555 2.825 0.555 2.825 0.54 2.945 0.54 2.945 0.555 3.265 0.555 3.265 0.495 3.325 0.495 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 1.19 1.66 1.19 1.66 0.93 1.5 0.93 1.5 0.85 1.74 0.85 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.92556625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.715 0.8 1.085 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.039375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.43809525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.02 0.925 0.96 0.925 0.96 1.245 0.475 1.245 0.475 1.11 0.26 1.11 0.26 0.955 0.535 0.955 0.535 1.185 0.9 1.185 0.9 0.865 1.02 0.865 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 1.77 0 1.77 0 1.65 0.605 1.65 0.605 1.345 0.725 1.345 0.725 1.405 0.665 1.405 0.665 1.65 1.76 1.65 1.76 1.29 1.82 1.29 1.82 1.65 2.24 1.65 2.24 1.15 2.3 1.15 2.3 1.65 2.65 1.65 2.65 1.15 2.71 1.15 2.71 1.65 3.06 1.65 3.06 1.15 3.12 1.15 3.12 1.65 3.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 0.06 3.12 0.06 3.12 0.455 3.06 0.455 3.06 0.06 2.71 0.06 2.71 0.455 2.65 0.455 2.65 0.06 2.295 0.06 2.295 0.455 2.235 0.455 2.235 0.06 1.635 0.06 1.635 0.365 1.695 0.365 1.695 0.425 1.575 0.425 1.575 0.06 0.695 0.06 0.695 0.455 0.635 0.455 0.635 0.06 0 0.06 0 -0.06 3.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.96 0.81 1.9 0.81 1.9 0.75 1.4 0.75 1.4 1.19 1.145 1.19 1.145 1.435 1.085 1.435 1.085 1.13 1.34 1.13 1.34 0.455 1.19 0.455 1.19 0.335 1.25 0.335 1.25 0.395 1.4 0.395 1.4 0.69 1.96 0.69 ;
      POLYGON 1.24 0.695 1.18 0.695 1.18 0.97 1.24 0.97 1.24 1.03 1.12 1.03 1.12 0.615 0.16 0.615 0.16 1.21 0.375 1.21 0.375 1.33 0.315 1.33 0.315 1.27 0.1 1.27 0.1 0.555 0.4 0.555 0.4 0.42 0.46 0.42 0.46 0.555 1.18 0.555 1.18 0.635 1.24 0.635 ;
  END
END MX2X8

MACRO MX2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX2XL 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6708 LAYER Metal1 ;
    ANTENNADIFFAREA 0.6762 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 20.70370375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 169.537037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.545 1.33 0.545 1.33 1.12 1.34 1.12 1.34 1.3 1.165 1.3 1.165 1.12 1.27 1.12 1.27 0.545 1.25 0.545 1.25 0.52 1.165 0.52 1.165 0.4 1.34 0.4 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.885 0.6 1.165 0.73 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.12962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.695 0.42 0.895 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.175926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.57 1.115 0.165 1.115 0.165 1.045 0.185 1.045 0.185 0.96 0.245 0.96 0.245 1.035 0.43 1.035 0.43 0.98 0.51 0.98 0.51 0.82 0.57 0.82 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.225 0.335 1.225 0.335 1.65 0.96 1.65 0.96 1.225 1.02 1.225 1.02 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 1.02 0.06 1.02 0.495 0.96 0.495 0.96 0.06 0.335 0.06 0.335 0.495 0.275 0.495 0.275 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.065 1.13 0.86 1.13 0.86 1.245 0.57 1.245 0.57 1.185 0.8 1.185 0.8 0.865 0.755 0.865 0.755 0.495 0.59 0.495 0.59 0.375 0.65 0.375 0.65 0.435 0.815 0.435 0.815 0.785 0.86 0.785 0.86 1.07 1.005 1.07 1.005 0.95 1.065 0.95 ;
      POLYGON 0.74 1.045 0.63 1.045 0.63 0.69 0.515 0.69 0.515 0.63 0.105 0.63 0.105 1.225 0.13 1.225 0.13 1.345 0.07 1.345 0.07 1.285 0.045 1.285 0.045 0.57 0.07 0.57 0.07 0.375 0.13 0.375 0.13 0.57 0.69 0.57 0.69 0.925 0.74 0.925 ;
  END
END MX2XL

MACRO MX3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX3X1 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4589 LAYER Metal1 ;
    ANTENNADIFFAREA 1.5071 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06165 LAYER Metal1 ;
      ANTENNAMAXAREACAR 23.6642335 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 187.88321175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.19 0.505 0.14 0.505 0.14 0.765 0.19 0.765 0.19 1.345 0.13 1.345 0.13 0.825 0.08 0.825 0.08 0.54 0.06 0.54 0.06 0.41 0.13 0.41 0.13 0.385 0.19 0.385 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.45370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.765 1.085 2.08 1.085 2.08 0.965 2.16 0.965 2.16 1.005 2.765 1.005 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.71 0.855 2.34 0.855 2.34 0.905 2.26 0.905 2.26 0.775 2.71 0.775 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.66 0.98 1.58 0.98 1.58 0.73 1.46 0.73 1.46 0.6 1.54 0.6 1.54 0.65 1.66 0.65 ;
    END
  END B
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.48 1.34 0.98 ;
    END
  END S1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.625 0.54 1.125 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.77 0 1.77 0 1.65 0.335 1.65 0.335 1.225 0.395 1.225 0.395 1.65 1.57 1.65 1.57 1.24 1.63 1.24 1.63 1.65 2.355 1.65 2.355 1.24 2.415 1.24 2.415 1.65 3 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 0.06 2.48 0.06 2.48 0.41 2.54 0.41 2.54 0.47 2.42 0.47 2.42 0.06 1.705 0.06 1.705 0.5 1.645 0.5 1.645 0.06 0.365 0.06 0.365 0.305 0.425 0.305 0.425 0.365 0.305 0.365 0.305 0.06 0 0.06 0 -0.06 3 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.925 1.245 2.66 1.245 2.66 1.305 2.6 1.305 2.6 1.185 2.865 1.185 2.865 0.675 2.16 0.675 2.16 0.82 1.98 0.82 1.98 0.975 1.92 0.975 1.92 0.76 2.1 0.76 2.1 0.615 2.865 0.615 2.865 0.515 2.655 0.515 2.655 0.395 2.715 0.395 2.715 0.455 2.925 0.455 ;
      POLYGON 2.23 0.495 2 0.495 2 0.66 1.82 0.66 1.82 1.08 1.98 1.08 1.98 1.185 2.045 1.185 2.045 1.305 1.985 1.305 1.985 1.245 1.92 1.245 1.92 1.14 1.055 1.14 1.055 0.32 1.175 0.32 1.175 0.38 1.115 0.38 1.115 1.08 1.76 1.08 1.76 0.6 1.94 0.6 1.94 0.435 2.23 0.435 ;
      POLYGON 1.5 0.5 1.44 0.5 1.44 0.22 0.955 0.22 0.955 1.3 1.365 1.3 1.365 1.24 1.425 1.24 1.425 1.36 0.895 1.36 0.895 0.89 0.835 0.89 0.835 0.77 0.895 0.77 0.895 0.595 0.835 0.595 0.835 0.535 0.895 0.535 0.895 0.16 1.5 0.16 ;
      POLYGON 0.795 0.405 0.735 0.405 0.735 0.99 0.795 0.99 0.795 1.05 0.675 1.05 0.675 0.525 0.36 0.525 0.36 0.665 0.24 0.665 0.24 0.605 0.3 0.605 0.3 0.465 0.675 0.465 0.675 0.345 0.795 0.345 ;
  END
END MX3X1

MACRO MX3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX3X2 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5441 LAYER Metal1 ;
    ANTENNADIFFAREA 1.743075 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0909 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.98679875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 134.37293725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.415 0.52 0.37 0.52 0.37 0.89 0.415 0.89 0.415 1.48 0.355 1.48 0.355 0.95 0.31 0.95 0.31 0.705 0.235 0.705 0.235 0.625 0.31 0.625 0.31 0.46 0.355 0.46 0.355 0.4 0.415 0.4 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.94 1.155 2.405 1.155 2.405 1.025 2.485 1.025 2.485 1.075 2.86 1.075 2.86 0.98 2.94 0.98 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.74 0.975 2.66 0.975 2.66 0.82 2.395 0.82 2.395 0.74 2.74 0.74 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.975 0.87 1.94 0.87 1.94 0.985 1.86 0.985 1.86 0.79 1.895 0.79 1.895 0.52 1.975 0.52 ;
    END
  END B
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.52 1.74 1.02 ;
    END
  END S1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.79 1.085 0.515 1.085 0.515 1.005 0.71 1.005 0.71 0.78 0.79 0.78 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 1.77 0 1.77 0 1.65 0.15 1.65 0.15 1.09 0.21 1.09 0.21 1.65 0.64 1.65 0.64 1.185 0.7 1.185 0.7 1.65 1.84 1.65 1.84 1.28 1.9 1.28 1.9 1.65 2.725 1.65 2.725 1.28 2.785 1.28 2.785 1.65 3.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 0.06 2.785 0.06 2.785 0.42 2.725 0.42 2.725 0.06 1.9 0.06 1.9 0.42 1.84 0.42 1.84 0.06 0.67 0.06 0.67 0.43 0.73 0.43 0.73 0.49 0.61 0.49 0.61 0.06 0.21 0.06 0.21 0.52 0.15 0.52 0.15 0.06 0 0.06 0 -0.06 3.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.1 1.315 2.995 1.315 2.995 1.375 2.935 1.375 2.935 1.255 3.04 1.255 3.04 0.64 2.295 0.64 2.295 1.02 2.235 1.02 2.235 0.58 2.49 0.58 2.49 0.52 2.55 0.52 2.55 0.58 3.04 0.58 3.04 0.445 2.935 0.445 2.935 0.325 2.995 0.325 2.995 0.385 3.1 0.385 ;
      POLYGON 2.475 0.42 2.135 0.42 2.135 1.255 2.37 1.255 2.37 1.375 2.31 1.375 2.31 1.315 2.075 1.315 2.075 1.18 1.37 1.18 1.37 1.12 1.475 1.12 1.475 0.63 1.405 0.63 1.405 0.57 1.535 0.57 1.535 1.12 2.075 1.12 2.075 0.36 2.415 0.36 2.415 0.3 2.475 0.3 ;
      POLYGON 1.725 1.34 1.21 1.34 1.21 0.95 1.11 0.95 1.11 1.01 1.05 1.01 1.05 0.89 1.315 0.89 1.315 0.79 1.245 0.79 1.245 0.3 1.695 0.3 1.695 0.42 1.635 0.42 1.635 0.36 1.305 0.36 1.305 0.73 1.375 0.73 1.375 0.95 1.27 0.95 1.27 1.28 1.725 1.28 ;
      POLYGON 1.145 0.68 0.95 0.68 0.95 1.11 1.105 1.11 1.105 1.23 1.045 1.23 1.045 1.17 0.89 1.17 0.89 0.68 0.59 0.68 0.59 0.79 0.47 0.79 0.47 0.62 1.085 0.62 1.085 0.54 1.145 0.54 ;
  END
END MX3X2

MACRO MX3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX3X4 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.87735 LAYER Metal1 ;
    ANTENNADIFFAREA 2.321525 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.16245 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.556479 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 88.531856 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.985 0.5 0.94 0.5 0.94 0.66 0.575 0.66 0.575 1.02 0.985 1.02 0.985 1.41 0.925 1.41 0.925 1.08 0.575 1.08 0.575 1.41 0.515 1.41 0.515 0.73 0.46 0.73 0.46 0.6 0.515 0.6 0.515 0.52 0.575 0.52 0.575 0.6 0.88 0.6 0.88 0.44 0.925 0.44 0.925 0.38 0.985 0.38 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.54 1.11 2.98 1.11 2.98 0.99 3.06 0.99 3.06 1.03 3.46 1.03 3.46 0.98 3.54 0.98 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.54 0.75 3.34 0.75 3.34 0.93 3.26 0.93 3.26 0.75 3.22 0.75 3.22 0.67 3.54 0.67 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.46 0.485 2.54 0.985 ;
    END
  END B
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.82838275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.485 2.34 0.985 ;
    END
  END S1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.41 0.84 1.34 0.84 1.34 1.19 1.26 1.19 1.26 0.76 1.41 0.76 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 1.77 0 1.77 0 1.65 0.3 1.65 0.3 1.02 0.36 1.02 0.36 1.65 0.72 1.65 0.72 1.18 0.78 1.18 0.78 1.65 1.21 1.65 1.21 1.29 1.27 1.29 1.27 1.65 2.41 1.65 2.41 1.245 2.47 1.245 2.47 1.65 3.295 1.65 3.295 1.275 3.415 1.275 3.415 1.335 3.355 1.335 3.355 1.65 3.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 0.06 3.385 0.06 3.385 0.385 3.325 0.385 3.325 0.06 2.475 0.06 2.475 0.385 2.415 0.385 2.415 0.06 1.27 0.06 1.27 0.5 1.21 0.5 1.21 0.06 0.78 0.06 0.78 0.5 0.72 0.5 0.72 0.06 0.37 0.06 0.37 0.5 0.31 0.5 0.31 0.06 0 0.06 0 -0.06 3.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.76 1.24 3.64 1.24 3.64 0.57 3.12 0.57 3.12 0.89 2.86 0.89 2.86 0.985 2.8 0.985 2.8 0.83 3.06 0.83 3.06 0.51 3.64 0.51 3.64 0.29 3.7 0.29 3.7 1.18 3.76 1.18 ;
      POLYGON 3.055 0.41 2.96 0.41 2.96 0.73 2.7 0.73 2.7 1.21 2.93 1.21 2.93 1.27 2.64 1.27 2.64 1.145 1.875 1.145 1.875 1.085 2.095 1.085 2.095 0.64 2.01 0.64 2.01 0.52 2.07 0.52 2.07 0.58 2.155 0.58 2.155 1.085 2.64 1.085 2.64 0.67 2.9 0.67 2.9 0.35 2.995 0.35 2.995 0.29 3.055 0.29 ;
      POLYGON 2.295 1.305 1.715 1.305 1.715 0.945 1.67 0.945 1.67 0.825 1.73 0.825 1.73 0.885 1.85 0.885 1.85 0.265 2.27 0.265 2.27 0.385 2.21 0.385 2.21 0.325 1.91 0.325 1.91 0.74 1.995 0.74 1.995 0.86 1.91 0.86 1.91 0.945 1.775 0.945 1.775 1.245 2.295 1.245 ;
      POLYGON 1.75 0.66 1.57 0.66 1.57 1.045 1.615 1.045 1.615 1.41 1.555 1.41 1.555 1.105 1.51 1.105 1.51 0.66 1.16 0.66 1.16 0.77 1.04 0.77 1.04 0.6 1.69 0.6 1.69 0.52 1.75 0.52 ;
  END
END MX3X4

MACRO MX3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX3XL 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.374975 LAYER Metal1 ;
    ANTENNADIFFAREA 1.437725 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXAREACAR 28.29166675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 225.2469135 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.16 1.29 0.04 1.29 0.04 1.23 0.1 1.23 0.1 0.54 0.06 0.54 0.06 0.41 0.16 0.41 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.7685185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.54 1.165 2.025 1.165 2.025 0.91 1.965 0.91 1.965 0.79 2.045 0.79 2.045 0.83 2.105 0.83 2.105 1.085 2.46 1.085 2.46 0.98 2.54 0.98 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.54 0.82 2.34 0.82 2.34 0.985 2.26 0.985 2.26 0.82 2.205 0.82 2.205 0.74 2.54 0.74 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.545 1.07 1.465 1.07 1.465 0.775 1.46 0.775 1.46 0.575 1.54 0.575 1.54 0.6 1.545 0.6 ;
    END
  END B
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 1.07 1.255 1.07 1.255 0.95 1.26 0.95 1.26 0.575 1.34 0.575 ;
    END
  END S1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.41 0.885 0.34 0.885 0.34 1.195 0.26 1.195 0.26 0.765 0.41 0.765 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 1.77 0 1.77 0 1.65 0.31 1.65 0.31 1.295 0.37 1.295 0.37 1.65 1.46 1.65 1.46 1.33 1.52 1.33 1.52 1.65 2.355 1.65 2.355 1.33 2.415 1.33 2.415 1.65 2.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 0.06 2.415 0.06 2.415 0.475 2.355 0.475 2.355 0.06 1.52 0.06 1.52 0.475 1.46 0.475 1.46 0.06 0.39 0.06 0.39 0.505 0.33 0.505 0.33 0.06 0 0.06 0 -0.06 2.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.7 1.355 2.64 1.355 2.64 0.64 2.105 0.64 2.105 0.69 1.865 0.69 1.865 1.01 1.925 1.01 1.925 1.07 1.805 1.07 1.805 0.63 1.985 0.63 1.985 0.595 2.06 0.595 2.06 0.58 2.64 0.58 2.64 0.38 2.7 0.38 ;
      POLYGON 1.995 0.495 1.705 0.495 1.705 1.235 1.945 1.235 1.945 1.355 1.885 1.355 1.885 1.295 1.645 1.295 1.645 1.23 1.155 1.23 1.155 1.29 0.99 1.29 0.99 1.23 1.095 1.23 1.095 0.53 1.055 0.53 1.055 0.41 1.115 0.41 1.115 0.47 1.155 0.47 1.155 1.17 1.645 1.17 1.645 0.435 1.935 0.435 1.935 0.375 1.995 0.375 ;
      POLYGON 1.315 0.475 1.255 0.475 1.255 0.31 0.955 0.31 0.955 0.63 0.995 0.63 0.995 0.75 0.955 0.75 0.955 1.07 0.89 1.07 0.89 1.39 1.255 1.39 1.255 1.33 1.315 1.33 1.315 1.45 0.83 1.45 0.83 1.07 0.73 1.07 0.73 1.13 0.67 1.13 0.67 1.01 0.895 1.01 0.895 0.25 1.315 0.25 ;
      POLYGON 0.795 0.665 0.57 0.665 0.57 1.23 0.73 1.23 0.73 1.29 0.51 1.29 0.51 0.665 0.26 0.665 0.26 0.605 0.735 0.605 0.735 0.41 0.795 0.41 ;
  END
END MX3XL

MACRO MX4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX4X1 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2257 LAYER Metal1 ;
    ANTENNADIFFAREA 2.224 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.07785 LAYER Metal1 ;
      ANTENNAMAXAREACAR 28.5895955 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 225.4913295 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.16 1.375 0.1 1.375 0.1 0.85 0.08 0.85 0.08 0.54 0.06 0.54 0.06 0.41 0.14 0.41 0.14 0.79 0.16 0.79 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.87654325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.165 0.895 3.565 0.895 3.565 1.405 2.405 1.405 2.405 1.345 3.505 1.345 3.505 0.905 3.445 0.905 3.445 0.835 4.035 0.835 4.035 0.815 4.165 0.815 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.935 0.735 3.615 0.735 3.615 0.705 3.465 0.705 3.465 0.625 3.765 0.625 3.765 0.655 3.935 0.655 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.135 1.085 2.835 1.085 2.835 1.005 2.885 1.005 2.885 0.805 2.965 0.805 2.965 1.005 3.135 1.005 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.735 1.085 2.435 1.085 2.435 1.005 2.655 1.005 2.655 0.805 2.735 0.805 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.015 1.01 1.885 1.01 1.885 0.705 1.82 0.705 1.82 0.625 1.965 0.625 1.965 0.835 2.015 0.835 ;
    END
  END D
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.625 0.98 0.505 0.98 0.505 0.705 0.4 0.705 0.4 0.625 0.565 0.625 0.565 0.645 0.625 0.645 ;
    END
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.305 1.65 0.305 1.08 0.365 1.08 0.365 1.65 1.895 1.65 1.895 1.27 1.955 1.27 1.955 1.65 2.755 1.65 2.755 1.54 2.875 1.54 2.875 1.65 3.72 1.65 3.72 1.07 3.78 1.07 3.78 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 3.79 0.06 3.79 0.365 3.67 0.365 3.67 0.305 3.73 0.305 3.73 0.06 2.875 0.06 2.875 0.525 2.815 0.525 2.815 0.06 2.195 0.06 2.195 0.305 2.255 0.305 2.255 0.365 2.135 0.365 2.135 0.06 0.335 0.06 0.335 0.305 0.395 0.305 0.395 0.365 0.275 0.365 0.275 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.325 1.055 3.995 1.055 3.995 1.115 3.935 1.115 3.935 0.995 4.265 0.995 4.265 0.525 3.51 0.525 3.51 0.25 3.125 0.25 3.125 0.76 3.185 0.76 3.185 0.82 3.065 0.82 3.065 0.705 2.335 0.705 2.335 0.85 2.275 0.85 2.275 0.645 3.065 0.645 3.065 0.19 3.57 0.19 3.57 0.465 3.935 0.465 3.935 0.405 3.995 0.405 3.995 0.465 4.325 0.465 ;
      POLYGON 3.345 1.245 2.055 1.245 2.055 1.17 1.6 1.17 1.6 0.8 1.66 0.8 1.66 0.54 1.535 0.54 1.535 0.42 1.595 0.42 1.595 0.48 1.72 0.48 1.72 0.86 1.66 0.86 1.66 1.11 2.115 1.11 2.115 1.185 3.285 1.185 3.285 0.52 3.225 0.52 3.225 0.46 3.345 0.46 ;
      POLYGON 2.565 0.525 2.175 0.525 2.175 0.95 2.275 0.95 2.275 1.005 2.335 1.005 2.335 1.065 2.215 1.065 2.215 1.01 2.115 1.01 2.115 0.525 1.975 0.525 1.975 0.32 1.18 0.32 1.18 0.99 1.045 0.99 1.045 0.93 1.12 0.93 1.12 0.26 2.035 0.26 2.035 0.465 2.505 0.465 2.505 0.405 2.565 0.405 ;
      POLYGON 1.56 0.7 1.5 0.7 1.5 1.33 0.665 1.33 0.665 1.08 0.725 1.08 0.725 0.505 0.655 0.505 0.655 0.445 0.785 0.445 0.785 1.14 0.725 1.14 0.725 1.27 1.44 1.27 1.44 0.64 1.56 0.64 ;
      POLYGON 1.385 0.545 1.34 0.545 1.34 1.15 0.885 1.15 0.885 0.345 0.555 0.345 0.555 0.525 0.3 0.525 0.3 0.72 0.24 0.72 0.24 0.465 0.495 0.465 0.495 0.285 0.945 0.285 0.945 1.09 1.28 1.09 1.28 0.485 1.325 0.485 1.325 0.425 1.385 0.425 ;
  END
END MX4X1

MACRO MX4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX4X2 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4841 LAYER Metal1 ;
    ANTENNADIFFAREA 2.871875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1071 LAYER Metal1 ;
      ANTENNAMAXAREACAR 23.194211 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 178.58543425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.75 0.68 1.74 0.68 1.74 1.04 1.6 1.04 1.6 0.96 1.66 0.96 1.66 0.6 1.67 0.6 1.67 0.425 1.75 0.425 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.099 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.037037 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 26.7901235 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.74 0.92 4.66 0.92 4.66 0.65 4.1 0.65 4.1 0.71 4.04 0.71 4.04 0.59 4.72 0.59 4.72 0.79 4.74 0.79 ;
    END
  END S0
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.56 0.895 4.28 0.895 4.28 0.97 4.2 0.97 4.2 0.75 4.56 0.75 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 1.06 3.34 1.06 3.34 1.28 3.26 1.28 3.26 0.98 3.32 0.98 3.32 0.84 3.4 0.84 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.28 2.86 1.28 2.86 0.965 2.92 0.965 2.92 0.84 3 0.84 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.175 0.87 1.94 0.87 1.94 0.92 1.86 0.92 1.86 0.79 2.095 0.79 2.095 0.655 2.175 0.655 ;
    END
  END A
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.73 1.27 0.73 1.27 0.87 1.17 0.87 1.17 0.62 1.26 0.62 1.26 0.46 1.34 0.46 ;
    END
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 1.77 0 1.77 0 1.65 1.365 1.65 1.365 1.54 1.485 1.54 1.485 1.65 1.835 1.65 1.835 1.3 1.955 1.3 1.955 1.36 1.895 1.36 1.895 1.65 3.015 1.65 3.015 1.54 3.135 1.54 3.135 1.65 4.285 1.65 4.285 1.23 4.345 1.23 4.345 1.65 5 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 0.06 4.315 0.06 4.315 0.43 4.375 0.43 4.375 0.49 4.255 0.49 4.255 0.06 3.2 0.06 3.2 0.36 3.08 0.36 3.08 0.3 3.14 0.3 3.14 0.06 2.07 0.06 2.07 0.2 2.01 0.2 2.01 0.06 1.41 0.06 1.41 0.2 1.35 0.2 1.35 0.06 0 0.06 0 -0.06 5 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.9 1.13 4.795 1.13 4.795 1.255 4.735 1.255 4.735 1.13 4.16 1.13 4.16 1.45 3.72 1.45 3.72 1.44 2.7 1.44 2.7 0.975 2.76 0.975 2.76 1.38 3.72 1.38 3.72 0.62 3.78 0.62 3.78 1.39 4.1 1.39 4.1 1.12 4.04 1.12 4.04 0.965 4.1 0.965 4.1 1.06 4.14 1.06 4.14 1.07 4.84 1.07 4.84 0.69 4.82 0.69 4.82 0.425 4.88 0.425 4.88 0.63 4.9 0.63 ;
      POLYGON 4 1.29 3.88 1.29 3.88 0.52 2.92 0.52 2.92 0.3 2.66 0.3 2.66 0.36 1.85 0.36 1.85 0.325 1.57 0.325 1.57 0.36 1.19 0.36 1.19 0.325 0.89 0.325 0.89 0.99 0.87 0.99 0.87 1.05 0.81 1.05 0.81 0.93 0.83 0.93 0.83 0.265 1.25 0.265 1.25 0.3 1.51 0.3 1.51 0.265 1.91 0.265 1.91 0.3 2.6 0.3 2.6 0.24 2.98 0.24 2.98 0.46 3.88 0.46 3.88 0.4 3.94 0.4 3.94 1.23 4 1.23 ;
      POLYGON 3.62 0.825 3.5 0.825 3.5 0.74 2.495 0.74 2.495 0.975 2.435 0.975 2.435 0.68 2.835 0.68 2.835 0.62 2.895 0.62 2.895 0.68 3.62 0.68 ;
      POLYGON 2.82 0.52 2.335 0.52 2.335 1.165 2.6 1.165 2.6 1.225 2.275 1.225 2.275 1.2 1.735 1.2 1.735 1.37 0.35 1.37 0.35 1.06 0.19 1.06 0.19 0.435 0.25 0.435 0.25 1 0.41 1 0.41 1.31 1.675 1.31 1.675 1.14 2.275 1.14 2.275 0.46 2.76 0.46 2.76 0.4 2.82 0.4 ;
      POLYGON 1.56 0.86 1.5 0.86 1.5 1.21 0.605 1.21 0.605 1.02 0.51 1.02 0.51 0.435 0.57 0.435 0.57 0.96 0.665 0.96 0.665 1.15 1.44 1.15 1.44 0.735 1.56 0.735 ;
      POLYGON 1.16 1.05 0.99 1.05 0.99 0.47 1.01 0.47 1.01 0.425 1.09 0.425 1.09 0.55 1.07 0.55 1.07 0.97 1.16 0.97 ;
      POLYGON 0.73 0.86 0.67 0.86 0.67 0.335 0.41 0.335 0.41 0.725 0.35 0.725 0.35 0.275 0.73 0.275 ;
  END
END MX4X2

MACRO MX4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX4X4 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0933 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.919753 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 25.771605 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.14 0.73 5.06 0.73 5.06 0.66 4.96 0.66 4.96 0.75 4.9 0.75 4.9 0.66 4.245 0.66 4.245 0.72 4.185 0.72 4.185 0.6 5.14 0.6 ;
    END
  END S0
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.895 4.485 0.895 4.485 1 4.405 1 4.405 0.815 4.8 0.815 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.765 1.085 3.465 1.085 3.465 0.805 3.545 0.805 3.545 1.005 3.765 1.005 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.14814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.235 0.805 3.365 1.115 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.46 0.53 2.54 1.03 ;
    END
  END A
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.82838275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.515 1.325 0.515 1.325 0.85 1.245 0.85 1.245 0.515 1.235 0.515 1.235 0.435 1.4 0.435 ;
    END
  END S1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7572 LAYER Metal1 ;
    ANTENNADIFFAREA 3.271825 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.17865 LAYER Metal1 ;
      ANTENNAMAXAREACAR 15.43352925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 117.74979 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.22 0.525 2.16 0.525 2.16 0.93 2.22 0.93 2.22 0.99 2.1 0.99 2.1 0.92 1.75 0.92 1.75 0.99 1.63 0.99 1.63 0.93 1.66 0.93 1.66 0.435 1.72 0.435 1.72 0.77 1.74 0.77 1.74 0.86 2.1 0.86 2.1 0.465 2.22 0.465 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 1.77 0 1.77 0 1.65 1.395 1.65 1.395 1.54 1.515 1.54 1.515 1.65 1.865 1.65 1.865 1.29 1.985 1.29 1.985 1.35 1.925 1.35 1.925 1.65 2.335 1.65 2.335 1.29 2.455 1.29 2.455 1.35 2.395 1.35 2.395 1.65 3.3 1.65 3.3 1.375 3.42 1.375 3.42 1.435 3.36 1.435 3.36 1.65 4.48 1.65 4.48 1.26 4.54 1.26 4.54 1.65 5.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 0.06 4.51 0.06 4.51 0.44 4.57 0.44 4.57 0.5 4.45 0.5 4.45 0.06 3.495 0.06 3.495 0.385 3.375 0.385 3.375 0.325 3.435 0.325 3.435 0.06 2.425 0.06 2.425 0.2 2.365 0.2 2.365 0.06 1.985 0.06 1.985 0.17 1.865 0.17 1.865 0.06 1.515 0.06 1.515 0.17 1.395 0.17 1.395 0.06 0 0.06 0 -0.06 5.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.3 1.16 5.035 1.16 5.035 1.285 4.975 1.285 4.975 1.16 4.305 1.16 4.305 1.415 3.865 1.415 3.865 1.275 3.065 1.275 3.065 1.04 3.025 1.04 3.025 0.92 3.085 0.92 3.085 0.97 3.125 0.97 3.125 1.215 3.865 1.215 3.865 0.645 3.925 0.645 3.925 1.355 4.245 1.355 4.245 1.085 4.185 1.085 4.185 1.025 4.305 1.025 4.305 1.1 5.24 1.1 5.24 0.5 4.945 0.5 4.945 0.44 5.3 0.44 ;
      POLYGON 4.145 1.255 4.025 1.255 4.025 0.545 3.215 0.545 3.215 0.325 2.955 0.325 2.955 0.36 2.205 0.36 2.205 0.335 0.895 0.335 0.895 0.95 0.955 0.95 0.955 1.01 0.835 1.01 0.835 0.275 2.265 0.275 2.265 0.3 2.895 0.3 2.895 0.265 3.275 0.265 3.275 0.485 4.025 0.485 4.025 0.425 4.085 0.425 4.085 1.195 4.145 1.195 ;
      POLYGON 3.765 0.85 3.645 0.85 3.645 0.705 2.86 0.705 2.86 1.005 2.8 1.005 2.8 0.645 3.765 0.645 ;
      POLYGON 3.115 0.545 2.7 0.545 2.7 1.13 2.965 1.13 2.965 1.255 2.845 1.255 2.845 1.19 1.765 1.19 1.765 1.35 0.355 1.35 0.355 0.96 0.195 0.96 0.195 0.43 0.255 0.43 0.255 0.9 0.415 0.9 0.415 1.29 1.705 1.29 1.705 1.13 2.64 1.13 2.64 0.485 3.055 0.485 3.055 0.425 3.115 0.425 ;
      POLYGON 1.56 0.85 1.485 0.85 1.485 1.19 0.635 1.19 0.635 1.01 0.515 1.01 0.515 0.43 0.575 0.43 0.575 0.95 0.695 0.95 0.695 1.13 1.425 1.13 1.425 0.79 1.5 0.79 1.5 0.73 1.56 0.73 ;
      POLYGON 1.28 1.03 1.055 1.03 1.055 0.85 0.995 0.85 0.995 0.73 1.055 0.73 1.055 0.435 1.135 0.435 1.135 0.95 1.28 0.95 ;
      POLYGON 0.735 0.85 0.675 0.85 0.675 0.33 0.415 0.33 0.415 0.715 0.355 0.715 0.355 0.27 0.735 0.27 ;
  END
END MX4X4

MACRO MX4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MX4XL 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1195 LAYER Metal1 ;
    ANTENNADIFFAREA 2.16495 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0648 LAYER Metal1 ;
      ANTENNAMAXAREACAR 32.70833325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 256.85185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.2 0.53 0.14 0.53 0.14 0.79 0.16 0.79 0.16 1.02 0.06 1.02 0.06 0.45 0.12 0.45 0.12 0.41 0.2 0.41 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.62962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.965 0.895 3.565 0.895 3.565 1.44 2.64 1.44 2.64 1.49 2.33 1.49 2.33 1.43 2.58 1.43 2.58 1.38 3.505 1.38 3.505 0.885 3.445 0.885 3.445 0.825 3.8 0.825 3.8 0.815 3.965 0.815 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.465 0.625 3.965 0.705 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.965 1.12 2.885 1.12 2.885 0.895 2.72 0.895 2.72 0.785 2.965 0.785 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.785 1.085 2.54 1.085 2.54 0.87 2.5 0.87 2.5 0.79 2.62 0.79 2.62 1.005 2.785 1.005 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.67 1.94 1.17 ;
    END
  END D
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 0.87 0.34 0.87 0.34 0.92 0.26 0.92 0.26 0.79 0.46 0.79 0.46 0.62 0.54 0.62 ;
    END
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 1.77 0 1.77 0 1.65 0.305 1.65 0.305 1.285 0.365 1.285 0.365 1.65 1.88 1.65 1.88 1.43 1.94 1.43 1.94 1.65 2.74 1.65 2.74 1.54 2.86 1.54 2.86 1.65 3.72 1.65 3.72 1.05 3.78 1.05 3.78 1.65 4.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 0.06 3.765 0.06 3.765 0.365 3.645 0.365 3.645 0.305 3.705 0.305 3.705 0.06 2.78 0.06 2.78 0.44 2.72 0.44 2.72 0.06 2.02 0.06 2.02 0.35 2.08 0.35 2.08 0.41 1.96 0.41 1.96 0.06 0.365 0.06 0.365 0.2 0.305 0.2 0.305 0.06 0 0.06 0 -0.06 4.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.125 1.11 4.02 1.11 4.02 1.17 3.96 1.17 3.96 1.05 4.065 1.05 4.065 0.525 3.445 0.525 3.445 0.23 3.125 0.23 3.125 0.705 3.185 0.705 3.185 0.765 3.065 0.765 3.065 0.685 2.4 0.685 2.4 0.73 2.26 0.73 2.26 0.84 2.2 0.84 2.2 0.67 2.34 0.67 2.34 0.625 3.065 0.625 3.065 0.17 3.505 0.17 3.505 0.465 3.91 0.465 3.91 0.345 3.97 0.345 3.97 0.465 4.125 0.465 ;
      POLYGON 3.345 1.015 3.23 1.015 3.23 1.28 2.48 1.28 2.48 1.33 1.515 1.33 1.515 0.54 1.575 0.54 1.575 1.27 2.42 1.27 2.42 1.22 3.17 1.22 3.17 0.955 3.285 0.955 3.285 0.435 3.225 0.435 3.225 0.375 3.345 0.375 ;
      POLYGON 2.47 0.465 2.24 0.465 2.24 0.57 2.1 0.57 2.1 0.94 2.26 0.94 2.26 0.985 2.32 0.985 2.32 1.045 2.2 1.045 2.2 1 2.04 1 2.04 0.57 1.675 0.57 1.675 0.44 1.05 0.44 1.05 1.02 1.08 1.02 1.08 1.08 0.96 1.08 0.96 1.02 0.99 1.02 0.99 0.38 1.735 0.38 1.735 0.51 2.18 0.51 2.18 0.405 2.41 0.405 2.41 0.345 2.47 0.345 ;
      POLYGON 1.415 1.425 0.64 1.425 0.64 0.43 0.7 0.43 0.7 1.365 1.355 1.365 1.355 0.7 1.415 0.7 ;
      POLYGON 1.255 1.24 0.8 1.24 0.8 0.33 0.525 0.33 0.525 0.52 0.36 0.52 0.36 0.69 0.24 0.69 0.24 0.63 0.3 0.63 0.3 0.46 0.465 0.46 0.465 0.27 0.86 0.27 0.86 1.18 1.195 1.18 1.195 0.54 1.255 0.54 ;
  END
END MX4XL

MACRO MXI2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X1 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6093 LAYER Metal1 ;
    ANTENNADIFFAREA 0.93715 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 20.83076925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 160.051282 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.855 0.545 0.72 0.545 0.72 0.79 0.74 0.79 0.74 0.92 0.72 0.92 0.72 1.365 0.66 1.365 0.66 0.485 0.855 0.485 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 12.87128725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 0.715 1.16 0.715 1.16 0.705 0.83 0.705 0.83 0.645 0.955 0.645 0.955 0.385 0.56 0.385 0.56 0.935 0.5 0.935 0.5 0.325 1.015 0.325 1.015 0.645 1.16 0.645 1.16 0.625 1.365 0.625 ;
    END
  END S0
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.41 0.895 1.14 0.895 1.14 0.985 1 0.985 1 0.815 1.41 0.815 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.535 0.34 1.035 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.255 1.65 0.255 1.135 0.315 1.135 0.315 1.65 1.085 1.65 1.085 1.245 1.145 1.245 1.145 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.175 0.06 1.175 0.525 1.115 0.525 1.115 0.06 0.315 0.06 0.315 0.435 0.255 0.435 0.255 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.57 1.145 1.35 1.145 1.35 1.27 1.29 1.27 1.29 1.145 0.84 1.145 0.84 0.815 0.9 0.815 0.9 1.085 1.51 1.085 1.51 0.525 1.32 0.525 1.32 0.405 1.38 0.405 1.38 0.465 1.57 0.465 ;
  END
END MXI2X1

MACRO MXI2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X2 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1561 LAYER Metal1 ;
    ANTENNADIFFAREA 1.44085 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0909 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.71837175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 95.8745875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 0.73 1.92 0.73 1.92 1.335 1.86 1.335 1.86 0.6 1.845 0.6 1.845 0.46 1.905 0.46 1.905 0.54 1.92 0.54 1.92 0.6 1.94 0.6 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.625 0.92 1.54 0.92 1.54 1.115 1.46 1.115 1.46 0.7 1.625 0.7 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.765 0.955 0.44 0.955 0.44 0.79 0.685 0.79 0.685 0.7 0.765 0.7 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.9 0.925 0.9 0.925 1.115 0.28 1.115 0.28 1.11 0.26 1.11 0.26 0.95 0.34 0.95 0.34 1.055 0.865 1.055 0.865 0.84 1.14 0.84 1.14 0.7 1.2 0.7 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 1.77 0 1.77 0 1.65 0.41 1.65 0.41 1.215 0.47 1.215 0.47 1.65 1.655 1.65 1.655 1.215 1.715 1.215 1.715 1.65 2.065 1.65 2.065 1.04 2.125 1.04 2.125 1.65 2.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 0.06 2.14 0.06 2.14 0.2 2.08 0.2 2.08 0.06 1.585 0.06 1.585 0.44 1.525 0.44 1.525 0.06 0.47 0.06 0.47 0.44 0.41 0.44 0.41 0.06 0 0.06 0 -0.06 2.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.405 0.55 2.345 0.55 2.345 0.675 2.375 0.675 2.375 1.065 2.315 1.065 2.315 0.735 2.04 0.735 2.04 0.675 2.285 0.675 2.285 0.49 2.405 0.49 ;
      POLYGON 2.36 0.355 2.3 0.355 2.3 0.36 1.745 0.36 1.745 0.6 1.36 0.6 1.36 1.06 1.085 1.06 1.085 1.24 1.025 1.24 1.025 1 1.3 1 1.3 0.46 1.075 0.46 1.075 0.34 1.135 0.34 1.135 0.4 1.36 0.4 1.36 0.54 1.685 0.54 1.685 0.3 2.24 0.3 2.24 0.295 2.36 0.295 ;
      POLYGON 1.005 0.66 0.945 0.66 0.945 0.6 0.16 0.6 0.16 1.215 0.265 1.215 0.265 1.335 0.205 1.335 0.205 1.275 0.1 1.275 0.1 0.54 0.205 0.54 0.205 0.345 0.265 0.345 0.265 0.54 1.005 0.54 ;
  END
END MXI2X2

MACRO MXI2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X4 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5005 LAYER Metal1 ;
    ANTENNADIFFAREA 1.828175 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.16245 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.23668825 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 71.44967675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.36 0.49 1.965 0.49 1.965 0.835 2.22 0.835 2.22 1.35 2.16 1.35 2.16 0.895 1.81 0.895 1.81 1.35 1.75 1.35 1.75 0.835 1.795 0.835 1.795 0.815 1.905 0.815 1.905 0.49 1.77 0.49 1.77 0.43 2.36 0.43 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 1.13 1.45 1.13 1.45 0.64 1.53 0.64 1.53 0.8 1.54 0.8 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.71 0.97 0.63 0.97 0.63 0.92 0.46 0.92 0.46 0.64 0.71 0.64 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 15.0925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.19 1.045 0.87 1.045 0.87 1.13 0.28 1.13 0.28 1.11 0.26 1.11 0.26 0.965 0.34 0.965 0.34 1.07 0.81 1.07 0.81 0.925 0.87 0.925 0.87 0.985 1.13 0.985 1.13 0.595 1.19 0.595 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.77 0 1.77 0 1.65 0.355 1.65 0.355 1.23 0.415 1.23 0.415 1.65 1.545 1.65 1.545 1.23 1.605 1.23 1.605 1.65 1.955 1.65 1.955 0.995 2.015 0.995 2.015 1.65 2.39 1.65 2.39 0.965 2.45 0.965 2.45 1.65 3 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 0.06 2.74 0.06 2.74 0.35 2.62 0.35 2.62 0.29 2.68 0.29 2.68 0.06 2.125 0.06 2.125 0.17 2.005 0.17 2.005 0.06 1.51 0.06 1.51 0.38 1.45 0.38 1.45 0.06 0.47 0.06 0.47 0.38 0.41 0.38 0.41 0.06 0 0.06 0 -0.06 3 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.915 0.52 2.75 0.52 2.75 0.865 2.655 0.865 2.655 1.35 2.595 1.35 2.595 0.865 2.32 0.865 2.32 0.805 2.69 0.805 2.69 0.46 2.855 0.46 2.855 0.4 2.915 0.4 ;
      POLYGON 2.59 0.705 2.53 0.705 2.53 0.51 2.46 0.51 2.46 0.33 1.67 0.33 1.67 0.54 1.35 0.54 1.35 1.29 0.955 1.29 0.955 1.35 0.895 1.35 0.895 1.23 1.29 1.23 1.29 0.38 1.065 0.38 1.065 0.26 1.125 0.26 1.125 0.32 1.35 0.32 1.35 0.48 1.61 0.48 1.61 0.27 2.52 0.27 2.52 0.45 2.59 0.45 ;
      POLYGON 1.03 0.885 0.97 0.885 0.97 0.54 0.16 0.54 0.16 1.18 0.18 1.18 0.18 1.3 0.12 1.3 0.12 1.23 0.1 1.23 0.1 0.48 0.205 0.48 0.205 0.285 0.265 0.285 0.265 0.48 1.03 0.48 ;
  END
END MXI2X4

MACRO MXI2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X6 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6484 LAYER Metal1 ;
    ANTENNADIFFAREA 2.008975 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2502 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.58832925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 52.18225425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.91 0.69 2.865 0.69 2.865 0.79 2.91 0.79 2.91 1.48 2.85 1.48 2.85 0.85 2.5 0.85 2.5 1.48 2.44 1.48 2.44 0.85 2.34 0.85 2.34 0.92 2.09 0.92 2.09 1.48 2.03 1.48 2.03 0.86 2.26 0.86 2.26 0.76 2.03 0.76 2.03 0.29 2.09 0.29 2.09 0.7 2.32 0.7 2.32 0.79 2.44 0.79 2.44 0.29 2.5 0.29 2.5 0.79 2.805 0.79 2.805 0.63 2.85 0.63 2.85 0.29 2.91 0.29 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.76 1.34 1.26 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.67 0.92 0.54 0.92 0.54 1.1 0.46 1.1 0.46 0.79 0.59 0.79 0.59 0.73 0.67 0.73 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.0925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.83 1.26 0.3 1.26 0.3 1.11 0.26 1.11 0.26 0.98 0.34 0.98 0.34 1.05 0.36 1.05 0.36 1.2 0.77 1.2 0.77 0.96 0.83 0.96 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.77 0 1.77 0 1.65 0.43 1.65 0.43 1.36 0.49 1.36 0.49 1.65 1.365 1.65 1.365 1.36 1.425 1.36 1.425 1.65 1.825 1.65 1.825 1.09 1.885 1.09 1.885 1.65 2.235 1.65 2.235 1.02 2.295 1.02 2.295 1.65 2.645 1.65 2.645 1.01 2.705 1.01 2.705 1.65 3 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 0.06 2.705 0.06 2.705 0.6 2.645 0.6 2.645 0.06 2.295 0.06 2.295 0.6 2.235 0.6 2.235 0.06 1.885 0.06 1.885 0.41 1.825 0.41 1.825 0.06 1.395 0.06 1.395 0.41 1.335 0.41 1.335 0.06 0.49 0.06 0.49 0.41 0.43 0.41 0.43 0.06 0 0.06 0 -0.06 3 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.93 0.76 1.725 0.76 1.725 1.15 1.63 1.15 1.63 1.48 1.57 1.48 1.57 1.09 1.665 1.09 1.665 0.5 1.57 0.5 1.57 0.38 1.63 0.38 1.63 0.44 1.725 0.44 1.725 0.7 1.93 0.7 ;
      POLYGON 1.565 0.72 1.505 0.72 1.505 0.66 1.16 0.66 1.16 1.355 0.93 1.355 0.93 1.295 1.1 1.295 1.1 0.41 0.8 0.41 0.8 0.29 0.86 0.29 0.86 0.35 1.16 0.35 1.16 0.6 1.565 0.6 ;
      POLYGON 1 1.195 0.94 1.195 0.94 0.82 0.93 0.82 0.93 0.63 0.16 0.63 0.16 1.2 0.2 1.2 0.2 1.385 0.14 1.385 0.14 1.26 0.1 1.26 0.1 0.375 0.225 0.375 0.225 0.315 0.285 0.315 0.285 0.435 0.16 0.435 0.16 0.57 0.76 0.57 0.76 0.51 0.99 0.51 0.99 0.76 1 0.76 ;
  END
END MXI2X6

MACRO MXI2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2X8 0 0 ;
  SIZE 3.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.825475 LAYER Metal1 ;
    ANTENNADIFFAREA 2.3541 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3078 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.930718 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 46.140351 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.35 0.51 2.97 0.51 2.97 0.98 3.35 0.98 3.35 1.425 3.29 1.425 3.29 1.04 2.94 1.04 2.94 1.425 2.88 1.425 2.88 1.04 2.53 1.04 2.53 1.425 2.47 1.425 2.47 1.04 2.14 1.04 2.14 1.11 2.12 1.11 2.12 1.425 2.06 1.425 2.06 0.405 2.12 0.405 2.12 0.98 2.91 0.98 2.91 0.51 2.515 0.51 2.515 0.495 2.44 0.495 2.44 0.435 2.56 0.435 2.56 0.45 2.85 0.45 2.85 0.435 2.97 0.435 2.97 0.45 3.29 0.45 3.29 0.39 3.35 0.39 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.705 1.34 1.205 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 0.92 0.54 0.92 0.54 1.025 0.46 1.025 0.46 0.645 0.66 0.645 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.861111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.84 1.205 0.28 1.205 0.28 1.11 0.26 1.11 0.26 0.98 0.34 0.98 0.34 0.99 0.36 0.99 0.36 1.125 0.76 1.125 0.76 0.865 0.84 0.865 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 1.77 0 1.77 0 1.65 0.43 1.65 0.43 1.305 0.49 1.305 0.49 1.65 1.395 1.65 1.395 1.305 1.455 1.305 1.455 1.65 1.855 1.65 1.855 1.035 1.915 1.035 1.915 1.65 2.265 1.65 2.265 1.14 2.325 1.14 2.325 1.65 2.675 1.65 2.675 1.14 2.735 1.14 2.735 1.65 3.085 1.65 3.085 1.14 3.145 1.14 3.145 1.65 3.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 0.06 3.145 0.06 3.145 0.35 3.085 0.35 3.085 0.06 2.735 0.06 2.735 0.35 2.675 0.35 2.675 0.06 2.325 0.06 2.325 0.35 2.265 0.35 2.265 0.06 1.915 0.06 1.915 0.385 1.855 0.385 1.855 0.06 1.395 0.06 1.395 0.385 1.335 0.385 1.335 0.06 0.49 0.06 0.49 0.385 0.43 0.385 0.43 0.06 0 0.06 0 -0.06 3.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.96 0.655 1.755 0.655 1.755 1.095 1.66 1.095 1.66 1.425 1.6 1.425 1.6 1.035 1.695 1.035 1.695 0.445 1.6 0.445 1.6 0.325 1.66 0.325 1.66 0.385 1.755 0.385 1.755 0.595 1.96 0.595 ;
      POLYGON 1.595 0.685 1.535 0.685 1.535 0.605 1.16 0.605 1.16 1.365 0.835 1.365 0.835 1.305 1.1 1.305 1.1 0.385 0.835 0.385 0.835 0.265 0.895 0.265 0.895 0.325 1.16 0.325 1.16 0.545 1.595 0.545 ;
      POLYGON 1 1.09 0.94 1.09 0.94 0.765 0.76 0.765 0.76 0.545 0.16 0.545 0.16 1.305 0.285 1.305 0.285 1.425 0.225 1.425 0.225 1.365 0.1 1.365 0.1 0.325 0.225 0.325 0.225 0.265 0.285 0.265 0.285 0.385 0.16 0.385 0.16 0.485 0.82 0.485 0.82 0.705 1 0.705 ;
  END
END MXI2X8

MACRO MXI2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI2XL 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5889 LAYER Metal1 ;
    ANTENNADIFFAREA 0.709675 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 36.35185175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 296.29629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.605 1.325 0.545 1.325 0.545 1.265 0.28 1.265 0.28 0.73 0.26 0.73 0.26 0.6 0.28 0.6 0.28 0.48 0.52 0.48 0.52 0.54 0.34 0.54 0.34 1.205 0.605 1.205 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.361111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.11 1.06 1.11 1.06 0.88 0.655 0.88 0.655 0.8 1.14 0.8 ;
    END
  END S0
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.77 0.98 0.96 1.2 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.18 1.2 0.1 1.2 0.1 0.92 0.06 0.92 0.06 0.74 0.14 0.74 0.14 0.84 0.18 0.84 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.12 1.65 0.12 1.3 0.18 1.3 0.18 1.65 0.93 1.65 0.93 1.3 0.99 1.3 0.99 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 0.96 0.06 0.96 0.48 1.02 0.48 1.02 0.54 0.9 0.54 0.9 0.06 0.22 0.06 0.22 0.2 0.16 0.2 0.16 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.3 1.325 1.24 1.325 1.24 0.7 0.555 0.7 0.555 0.98 0.67 0.98 0.67 1.1 0.61 1.1 0.61 1.04 0.495 1.04 0.495 0.64 0.62 0.64 0.62 0.38 0.385 0.38 0.385 0.27 0.325 0.27 0.325 0.21 0.445 0.21 0.445 0.32 0.68 0.32 0.68 0.64 1.135 0.64 1.135 0.475 1.195 0.475 1.195 0.64 1.3 0.64 ;
  END
END MXI2XL

MACRO MXI3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI3X1 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8423 LAYER Metal1 ;
    ANTENNADIFFAREA 2.028625 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.09405 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.58851675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 152.7910685 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.54 3.74 1.29 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 0.74 3.315 0.74 3.315 0.86 3.235 0.86 3.235 0.74 3.06 0.74 3.06 0.62 3.4 0.62 ;
    END
  END C
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.765 0.99 2.235 0.99 2.235 0.8 2.355 0.8 2.355 0.815 2.365 0.815 2.365 0.91 2.765 0.91 ;
    END
  END S1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.755 1.085 1.42 1.085 1.42 0.84 1.5 0.84 1.5 1.005 1.755 1.005 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.82 0.855 0.565 0.855 0.565 0.905 0.37 0.905 0.37 0.775 0.82 0.775 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.95370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.085 0.19 1.085 0.19 0.895 0.27 0.895 0.27 1.005 0.92 1.005 0.92 0.93 1 0.93 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 1.77 0 1.77 0 1.65 0.34 1.65 0.34 1.185 0.4 1.185 0.4 1.65 1.485 1.65 1.485 1.185 1.545 1.185 1.545 1.65 2.375 1.65 2.375 1.54 2.495 1.54 2.495 1.65 3.395 1.65 3.395 1.345 3.515 1.345 3.515 1.405 3.455 1.405 3.455 1.65 3.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 0.06 3.51 0.06 3.51 0.52 3.45 0.52 3.45 0.06 2.565 0.06 2.565 0.43 2.625 0.43 2.625 0.49 2.505 0.49 2.505 0.06 1.545 0.06 1.545 0.52 1.485 0.52 1.485 0.06 0.37 0.06 0.37 0.43 0.43 0.43 0.43 0.49 0.31 0.49 0.31 0.06 0 0.06 0 -0.06 3.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.56 1.02 3.41 1.02 3.41 1.245 3.295 1.245 3.295 1.34 1.915 1.34 1.915 1.18 1.855 1.18 1.855 0.455 1.975 0.455 1.975 0.515 1.915 0.515 1.915 1.12 1.975 1.12 1.975 1.28 3.235 1.28 3.235 1.185 3.35 1.185 3.35 0.96 3.5 0.96 3.5 0.74 3.56 0.74 ;
      POLYGON 3.305 0.52 2.96 0.52 2.96 1.025 3.25 1.025 3.25 1.085 2.9 1.085 2.9 0.81 2.465 0.81 2.465 0.75 2.9 0.75 2.9 0.46 3.245 0.46 3.245 0.4 3.305 0.4 ;
      POLYGON 2.8 0.65 2.345 0.65 2.345 0.355 2.135 0.355 2.135 1.12 2.73 1.12 2.73 1.18 2.075 1.18 2.075 1.02 2.015 1.02 2.015 0.96 2.075 0.96 2.075 0.355 1.85 0.355 1.85 0.26 1.79 0.26 1.79 0.2 1.91 0.2 1.91 0.295 2.405 0.295 2.405 0.59 2.74 0.59 2.74 0.425 2.8 0.425 ;
      POLYGON 1.62 0.74 1.32 0.74 1.32 1.245 1.03 1.245 1.03 1.185 1.26 1.185 1.26 0.515 0.825 0.515 0.825 0.455 1.32 0.455 1.32 0.68 1.56 0.68 1.56 0.62 1.62 0.62 ;
      POLYGON 1.16 0.965 1.1 0.965 1.1 0.675 0.09 0.675 0.09 1.185 0.195 1.185 0.195 1.305 0.135 1.305 0.135 1.245 0.03 1.245 0.03 0.615 0.135 0.615 0.135 0.425 0.195 0.425 0.195 0.615 1.16 0.615 ;
  END
END MXI3X1

MACRO MXI3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI3X2 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.669975 LAYER Metal1 ;
    ANTENNADIFFAREA 2.21195 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1233 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.5439985 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 102.1776155 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.17 0.65 2.14 0.65 2.14 1.335 2.06 1.335 2.06 0.65 2.05 0.65 2.05 0.57 2.17 0.57 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 15.60185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.565 0.705 3.435 0.705 3.435 0.55 2.96 0.55 2.96 0.68 2.9 0.68 2.9 0.55 2.75 0.55 2.75 0.9 2.695 0.9 2.695 0.96 2.635 0.96 2.635 0.84 2.69 0.84 2.69 0.49 3.555 0.49 3.555 0.625 3.565 0.625 ;
    END
  END S0
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.335 0.955 3.06 0.955 3.06 0.79 3.255 0.79 3.255 0.65 3.335 0.65 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.375 0.87 2.34 0.87 2.34 0.92 2.26 0.92 2.26 0.79 2.295 0.79 2.295 0.455 2.375 0.455 ;
    END
  END A
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.545 1.065 0.965 1.065 0.965 1.085 0.835 1.085 0.835 1.065 0.72 1.065 0.72 0.88 0.78 0.88 0.78 1.005 1.22 1.005 1.22 0.71 1.28 0.71 1.28 1.005 1.485 1.005 1.485 0.87 1.545 0.87 ;
    END
  END S1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.26 1.06 0.14 1.06 0.14 1.11 0.06 1.11 0.06 0.98 0.18 0.98 0.18 0.73 0.26 0.73 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 1.77 0 1.77 0 1.65 0.135 1.65 0.135 1.21 0.195 1.21 0.195 1.65 0.795 1.65 0.795 1.51 0.855 1.51 0.855 1.65 1.875 1.65 1.875 1.04 1.935 1.04 1.935 1.65 2.285 1.65 2.285 1.02 2.345 1.02 2.345 1.65 3.18 1.65 3.18 1.215 3.24 1.215 3.24 1.65 3.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 0.06 3.24 0.06 3.24 0.39 3.18 0.39 3.18 0.06 2.405 0.06 2.405 0.17 2.285 0.17 2.285 0.06 1.935 0.06 1.935 0.17 1.815 0.17 1.815 0.06 0.855 0.06 0.855 0.2 0.795 0.2 0.795 0.06 0.15 0.06 0.15 0.63 0.09 0.63 0.09 0.06 0 0.06 0 -0.06 3.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.725 1.115 3.445 1.115 3.445 1.24 3.385 1.24 3.385 1.115 2.85 1.115 2.85 0.96 2.91 0.96 2.91 1.055 3.665 1.055 3.665 0.39 3.54 0.39 3.54 0.27 3.6 0.27 3.6 0.33 3.725 0.33 ;
      POLYGON 2.93 0.39 2.87 0.39 2.87 0.33 2.535 0.33 2.535 1.215 2.8 1.215 2.8 1.275 2.475 1.275 2.475 0.33 1.595 0.33 1.595 0.27 2.93 0.27 ;
      POLYGON 1.96 0.83 1.9 0.83 1.9 0.77 1.705 0.77 1.705 1.225 1.38 1.225 1.38 1.165 1.645 1.165 1.645 0.77 1.38 0.77 1.38 0.54 1.44 0.54 1.44 0.71 1.96 0.71 ;
      POLYGON 1.12 0.905 1.06 0.905 1.06 0.78 0.62 0.78 0.62 1.16 0.56 1.16 0.56 0.54 0.62 0.54 0.62 0.72 1.12 0.72 ;
      POLYGON 1.075 0.445 0.82 0.445 0.82 0.44 0.42 0.44 0.42 1.235 0.36 1.235 0.36 0.38 0.855 0.38 0.855 0.385 1.075 0.385 ;
  END
END MXI3X2

MACRO MXI3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI3X4 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9811 LAYER Metal1 ;
    ANTENNADIFFAREA 2.444 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.202725 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.77235175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 75.10173875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.61 0.53 2.485 0.53 2.485 1.35 2.425 1.35 2.425 0.92 2.12 0.92 2.12 1.025 2.075 1.025 2.075 1.35 2.015 1.35 2.015 0.965 2.06 0.965 2.06 0.79 2.14 0.79 2.14 0.86 2.425 0.86 2.425 0.53 2.02 0.53 2.02 0.47 2.61 0.47 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.71 0.705 3.325 0.705 3.325 0.765 3.235 0.765 3.235 0.705 3.06 0.705 3.06 1.015 3 1.015 3 0.645 3.235 0.645 3.235 0.625 3.365 0.625 3.365 0.645 3.71 0.645 ;
    END
  END S0
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.77 0.945 3.33 0.945 3.33 0.865 3.635 0.865 3.635 0.805 3.77 0.805 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.66 0.63 2.74 1.13 ;
    END
  END A
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.039375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.14285725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.47 0.955 1.35 0.955 1.35 0.77 1.09 0.77 1.09 0.83 0.825 0.83 0.825 0.85 0.705 0.85 0.705 0.79 0.765 0.79 0.765 0.77 1.03 0.77 1.03 0.685 1.06 0.685 1.06 0.6 1.14 0.6 1.14 0.71 1.41 0.71 1.41 0.895 1.47 0.895 ;
    END
  END S1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.255 0.795 0.175 0.795 0.175 0.54 0.06 0.54 0.06 0.41 0.14 0.41 0.14 0.46 0.255 0.46 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 0 1.77 0 1.65 0.15 1.65 0.15 0.995 0.21 0.995 0.21 1.65 0.895 1.65 0.895 1.23 0.955 1.23 0.955 1.65 1.73 1.65 1.73 0.965 1.79 0.965 1.79 1.65 2.22 1.65 2.22 1.02 2.28 1.02 2.28 1.65 2.63 1.65 2.63 1.23 2.69 1.23 2.69 1.65 3.49 1.65 3.49 1.205 3.55 1.205 3.55 1.65 4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.605 0.06 3.605 0.525 3.545 0.525 3.545 0.06 2.845 0.06 2.845 0.17 2.725 0.17 2.725 0.06 2.375 0.06 2.375 0.17 2.255 0.17 2.255 0.06 1.76 0.06 1.76 0.42 1.7 0.42 1.7 0.06 0.965 0.06 0.965 0.42 0.905 0.42 0.905 0.06 0.25 0.06 0.25 0.2 0.19 0.2 0.19 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.93 1.105 3.755 1.105 3.755 1.23 3.695 1.23 3.695 1.105 3.17 1.105 3.17 0.95 3.23 0.95 3.23 1.045 3.87 1.045 3.87 0.43 3.93 0.43 ;
      POLYGON 3.295 0.525 3.235 0.525 3.235 0.465 2.9 0.465 2.9 1.115 3.07 1.115 3.07 1.235 3.01 1.235 3.01 1.175 2.84 1.175 2.84 0.465 2.71 0.465 2.71 0.37 1.92 0.37 1.92 0.635 1.67 0.635 1.67 0.575 1.86 0.575 1.86 0.31 2.77 0.31 2.77 0.405 3.295 0.405 ;
      POLYGON 1.96 0.865 1.63 0.865 1.63 1.15 1.365 1.15 1.365 1.35 1.305 1.35 1.305 1.09 1.57 1.09 1.57 0.795 1.51 0.795 1.51 0.61 1.24 0.61 1.24 0.385 1.3 0.385 1.3 0.55 1.57 0.55 1.57 0.735 1.63 0.735 1.63 0.805 1.96 0.805 ;
      POLYGON 1.25 0.99 0.985 0.99 0.985 1.01 0.72 1.01 0.72 1.16 0.66 1.16 0.66 1.01 0.525 1.01 0.525 0.415 0.645 0.415 0.645 0.475 0.585 0.475 0.585 0.95 0.925 0.95 0.925 0.93 1.19 0.93 1.19 0.87 1.25 0.87 ;
      POLYGON 0.93 0.67 0.745 0.67 0.745 0.315 0.415 0.315 0.415 1.02 0.355 1.02 0.355 0.255 0.805 0.255 0.805 0.61 0.93 0.61 ;
  END
END MXI3X4

MACRO MXI3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI3XL 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6611 LAYER Metal1 ;
    ANTENNADIFFAREA 1.736525 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.081 LAYER Metal1 ;
      ANTENNAMAXAREACAR 20.5074075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 160.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.52 3.34 1.02 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.15 1.085 2.915 1.085 2.915 0.74 2.995 0.74 2.995 0.79 3.15 0.79 ;
    END
  END C
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.8055555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.565 1.02 2.035 1.02 2.035 0.815 2.165 0.815 2.165 0.94 2.565 0.94 ;
    END
  END S1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.9814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.345 0.845 1.54 1.135 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.425 0.815 0.925 0.895 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.2685185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.9 1.075 0.365 1.075 0.365 1.085 0.235 1.085 0.235 1.005 0.245 1.005 0.245 0.965 0.325 0.965 0.325 0.995 0.9 0.995 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 1.77 0 1.77 0 1.65 0.5 1.65 0.5 1.235 0.56 1.235 0.56 1.65 1.375 1.65 1.375 1.235 1.435 1.235 1.435 1.65 2.175 1.65 2.175 1.54 2.295 1.54 2.295 1.65 2.995 1.65 2.995 1.345 3.115 1.345 3.115 1.405 3.055 1.405 3.055 1.65 3.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 0.06 3.115 0.06 3.115 0.635 3.055 0.635 3.055 0.06 2.365 0.06 2.365 0.46 2.425 0.46 2.425 0.52 2.305 0.52 2.305 0.06 1.405 0.06 1.405 0.46 1.465 0.46 1.465 0.52 1.345 0.52 1.345 0.06 0.56 0.06 0.56 0.55 0.5 0.55 0.5 0.06 0 0.06 0 -0.06 3.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.285 1.245 2.895 1.245 2.895 1.39 1.715 1.39 1.715 1.23 1.655 1.23 1.655 0.485 1.775 0.485 1.775 0.545 1.715 0.545 1.715 1.17 1.775 1.17 1.775 1.33 2.835 1.33 2.835 1.185 3.285 1.185 ;
      POLYGON 2.91 0.64 2.815 0.64 2.815 1.02 2.755 1.02 2.755 0.84 2.265 0.84 2.265 0.78 2.755 0.78 2.755 0.58 2.85 0.58 2.85 0.52 2.91 0.52 ;
      POLYGON 2.6 0.68 1.935 0.68 1.935 1.17 2.53 1.17 2.53 1.23 1.875 1.23 1.875 1.07 1.815 1.07 1.815 1.01 1.875 1.01 1.875 0.385 1.64 0.385 1.64 0.3 1.58 0.3 1.58 0.24 1.7 0.24 1.7 0.325 1.935 0.325 1.935 0.62 2.54 0.62 2.54 0.455 2.6 0.455 ;
      POLYGON 1.51 0.745 1.245 0.745 1.245 1.235 0.92 1.235 0.92 1.175 1.185 1.175 1.185 0.545 0.78 0.545 0.78 0.485 1.245 0.485 1.245 0.685 1.45 0.685 1.45 0.625 1.51 0.625 ;
      POLYGON 1.085 0.98 1.025 0.98 1.025 0.715 0.135 0.715 0.135 1.185 0.355 1.185 0.355 1.305 0.295 1.305 0.295 1.245 0.075 1.245 0.075 0.655 0.295 0.655 0.295 0.455 0.355 0.455 0.355 0.655 1.085 0.655 ;
  END
END MXI3XL

MACRO MXI4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI4X1 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.072 LAYER Metal1 ;
    ANTENNADIFFAREA 2.4234 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.11025 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.79365075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 141.904762 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.21 1.34 0.13 1.34 0.13 0.73 0.06 0.73 0.06 0.6 0.13 0.6 0.13 0.54 0.21 0.54 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0758 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.55967075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 15.43209875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.405 0.815 3.905 0.895 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.79 1.19 3.405 1.19 3.405 0.995 3.565 0.995 3.565 1.065 3.79 1.065 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.805 0.94 2.965 1.19 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.705 1.085 2.405 1.085 2.405 1.005 2.585 1.005 2.585 0.805 2.705 0.805 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.985 1 1.685 1 1.685 0.895 1.59 0.895 1.59 0.815 1.765 0.815 1.765 0.9 1.985 0.9 ;
    END
  END D
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 20.27777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.49 0.88 1.43 0.88 1.43 0.305 1.095 0.305 1.095 0.33 0.54 0.33 0.54 0.83 0.48 0.83 0.48 0.54 0.46 0.54 0.46 0.41 0.48 0.41 0.48 0.27 1.035 0.27 1.035 0.245 1.49 0.245 ;
    END
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 1.77 0 1.77 0 1.65 0.325 1.65 0.325 1.25 0.445 1.25 0.445 1.31 0.385 1.31 0.385 1.65 0.755 1.65 0.755 1.25 0.875 1.25 0.875 1.31 0.815 1.31 0.815 1.65 1.79 1.65 1.79 1.54 1.91 1.54 1.91 1.65 2.77 1.65 2.77 1.51 2.71 1.51 2.71 1.45 2.83 1.45 2.83 1.65 3.605 1.65 3.605 1.29 3.665 1.29 3.665 1.65 4.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 0.06 3.77 0.06 3.77 0.2 3.71 0.2 3.71 0.06 2.805 0.06 2.805 0.365 2.745 0.365 2.745 0.06 1.725 0.06 1.725 0.555 1.665 0.555 1.665 0.06 0.96 0.06 0.96 0.17 0.84 0.17 0.84 0.06 0.475 0.06 0.475 0.17 0.355 0.17 0.355 0.06 0 0.06 0 -0.06 4.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.065 1.255 3.95 1.255 3.95 1.315 3.89 1.315 3.89 1.195 4.005 1.195 4.005 0.36 3.465 0.36 3.465 0.23 3.145 0.23 3.145 1.045 3.085 1.045 3.085 0.525 2.585 0.525 2.585 0.22 2.145 0.22 2.145 0.985 2.085 0.985 2.085 0.16 2.645 0.16 2.645 0.465 3.085 0.465 3.085 0.17 3.525 0.17 3.525 0.3 4.065 0.3 ;
      POLYGON 3.365 0.55 3.305 0.55 3.305 1.41 3.245 1.41 3.245 1.35 2.465 1.35 2.465 1.44 1.57 1.44 1.57 1.38 2.405 1.38 2.405 1.29 3.245 1.29 3.245 0.49 3.365 0.49 ;
      POLYGON 2.985 0.84 2.865 0.84 2.865 0.705 2.485 0.705 2.485 0.87 2.405 0.87 2.405 0.625 2.985 0.625 ;
      POLYGON 2.44 0.525 2.305 0.525 2.305 1.22 2.245 1.22 2.245 1.16 1.53 1.16 1.53 1.28 1.47 1.28 1.47 1.37 1.095 1.37 1.095 1.375 0.975 1.375 0.975 1.315 1.035 1.315 1.035 1.31 1.41 1.31 1.41 1.22 1.47 1.22 1.47 1.1 2.245 1.1 2.245 0.465 2.44 0.465 ;
      POLYGON 1.33 1.12 1.31 1.12 1.31 1.21 1.25 1.21 1.25 1.15 0.31 1.15 0.31 0.74 0.37 0.74 0.37 1.09 1.25 1.09 1.25 1.06 1.27 1.06 1.27 0.55 1.18 0.55 1.18 0.49 1.33 0.49 ;
      POLYGON 1.17 0.99 0.58 0.99 0.58 0.93 0.7 0.93 0.7 0.63 0.64 0.63 0.64 0.57 0.76 0.57 0.76 0.93 1.11 0.93 1.11 0.87 1.17 0.87 ;
  END
END MXI4X1

MACRO MXI4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI4X2 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.63545 LAYER Metal1 ;
    ANTENNADIFFAREA 3.30585 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1395 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.89211475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 142.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.74 0.92 4.725 0.92 4.725 1.025 4.645 1.025 4.645 0.645 4.605 0.645 4.605 0.565 4.725 0.565 4.725 0.79 4.74 0.79 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.585 1.005 1.92 1.25 ;
    END
  END C
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0912 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.87654325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 24.87654325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.73 0.86 0.65 0.86 0.65 0.73 0.345 0.73 0.345 0.92 0.26 0.92 0.26 0.65 0.73 0.65 ;
    END
  END S0
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.485 1.25 1.15 1.25 1.15 1.005 1.365 1.005 1.365 1.015 1.485 1.015 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.73 1.04 0.54 1.04 0.54 1.14 0.46 1.14 0.46 0.83 0.54 0.83 0.54 0.96 0.73 0.96 ;
    END
  END A
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 27.4074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.165 0.895 5.02 0.895 5.02 1.315 3.305 1.315 3.305 0.875 3.39 0.875 3.39 0.79 3.45 0.79 3.45 0.935 3.365 0.935 3.365 1.255 4.96 1.255 4.96 0.835 5.035 0.835 5.035 0.765 5.165 0.765 ;
    END
  END S1
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.86 0.62 2.94 1.12 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 1.77 0 1.77 0 1.65 0.425 1.65 0.425 1.24 0.485 1.24 0.485 1.65 1.35 1.65 1.35 1.51 1.41 1.51 1.41 1.65 2.935 1.65 2.935 1.54 3.055 1.54 3.055 1.65 4.41 1.65 4.41 1.51 4.47 1.51 4.47 1.65 4.985 1.65 4.985 1.51 5.045 1.51 5.045 1.65 5.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 0.06 5.045 0.06 5.045 0.5 4.985 0.5 4.985 0.06 4.165 0.06 4.165 0.43 4.225 0.43 4.225 0.49 4.105 0.49 4.105 0.06 3.025 0.06 3.025 0.36 2.965 0.36 2.965 0.06 1.485 0.06 1.485 0.2 1.425 0.2 1.425 0.06 0.455 0.06 0.455 0.39 0.395 0.39 0.395 0.06 0 0.06 0 -0.06 5.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.325 1.055 5.12 1.055 5.12 0.995 5.265 0.995 5.265 0.66 4.825 0.66 4.825 0.465 4.385 0.465 4.385 0.995 3.625 0.995 3.625 0.69 3.285 0.69 3.285 0.63 3.685 0.63 3.685 0.935 4.325 0.935 4.325 0.405 4.885 0.405 4.885 0.6 5.22 0.6 5.22 0.54 5.325 0.54 ;
      POLYGON 4.545 1.155 3.465 1.155 3.465 1.035 3.525 1.035 3.525 1.095 4.485 1.095 4.485 0.745 4.545 0.745 ;
      POLYGON 4.225 0.835 3.785 0.835 3.785 0.53 3.415 0.53 3.415 0.515 3.355 0.515 3.355 0.455 3.475 0.455 3.475 0.47 3.845 0.47 3.845 0.775 4.225 0.775 ;
      POLYGON 4.065 0.675 3.945 0.675 3.945 0.355 3.185 0.355 3.185 0.52 2.76 0.52 2.76 1.28 2.415 1.28 2.415 1.22 2.7 1.22 2.7 0.52 2.325 0.52 2.325 0.4 2.385 0.4 2.385 0.46 3.125 0.46 3.125 0.295 4.005 0.295 4.005 0.615 4.065 0.615 ;
      POLYGON 3.185 1.44 1.51 1.44 1.51 1.41 0.83 1.41 0.83 0.425 0.89 0.425 0.89 1.35 1.57 1.35 1.57 1.38 3.125 1.38 3.125 0.79 3.185 0.79 ;
      POLYGON 2.6 1.12 2.48 1.12 2.48 1.04 2.18 1.04 2.18 0.96 2.56 0.96 2.56 1.015 2.6 1.015 ;
      POLYGON 2.48 0.855 2.4 0.855 2.4 0.86 2.08 0.86 2.08 0.985 2.02 0.985 2.02 0.86 1.15 0.86 1.15 0.74 1.21 0.74 1.21 0.8 2.34 0.8 2.34 0.795 2.48 0.795 ;
      RECT 1.74 0.62 2.24 0.7 ;
      POLYGON 1.86 0.28 1.645 0.28 1.645 0.36 1.265 0.36 1.265 0.325 1.05 0.325 1.05 1.02 0.99 1.02 0.99 0.325 0.7 0.325 0.7 0.55 0.16 0.55 0.16 1.02 0.28 1.02 0.28 1.265 0.22 1.265 0.22 1.08 0.1 1.08 0.1 0.49 0.16 0.49 0.16 0.43 0.22 0.43 0.22 0.49 0.64 0.49 0.64 0.16 0.76 0.16 0.76 0.265 1.325 0.265 1.325 0.3 1.585 0.3 1.585 0.22 1.86 0.22 ;
  END
END MXI4X2

MACRO MXI4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI4X4 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.039375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 26.05714275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.205 0.875 4.965 0.875 4.965 1.155 4.685 1.155 4.685 1.315 2.835 1.315 2.835 0.775 2.895 0.775 2.895 1.255 4.625 1.255 4.625 1.095 4.905 1.095 4.905 0.895 4.835 0.895 4.835 0.815 5.205 0.815 ;
    END
  END S1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8319 LAYER Metal1 ;
    ANTENNADIFFAREA 3.517575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.218925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.93548025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 99.7464885 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.84 0.645 4.54 0.645 4.54 0.935 4.67 0.935 4.67 0.995 4.48 0.995 4.48 0.73 4.46 0.73 4.46 0.645 4.2 0.645 4.2 0.995 4.08 0.995 4.08 0.935 4.14 0.935 4.14 0.645 4.08 0.645 4.08 0.375 4.14 0.375 4.14 0.585 4.78 0.585 4.78 0.375 4.84 0.375 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.575 1.2 2.46 1.2 2.46 1.1 2.445 1.1 2.445 0.75 2.525 0.75 2.525 0.98 2.575 0.98 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.76 1.2 1.66 1.2 1.66 0.98 1.68 0.98 1.68 0.72 1.76 0.72 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.56 1.1 1.54 1.1 1.54 1.2 1.46 1.2 1.46 0.98 1.48 0.98 1.48 0.72 1.56 0.72 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.865 0.58 1.205 ;
    END
  END A
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0843 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.734568 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 24.50617275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.89 0.94 0.81 0.94 0.81 0.765 0.34 0.765 0.34 0.92 0.26 0.92 0.26 0.685 0.89 0.685 ;
    END
  END S0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 0 1.77 0 1.65 0.41 1.65 0.41 1.305 0.47 1.305 0.47 1.65 1.47 1.65 1.47 1.46 1.59 1.46 1.59 1.52 1.53 1.52 1.53 1.65 2.51 1.65 2.51 1.46 2.63 1.46 2.63 1.52 2.57 1.52 2.57 1.65 3.645 1.65 3.645 1.54 3.765 1.54 3.765 1.65 4.315 1.65 4.315 1.54 4.435 1.54 4.435 1.65 4.785 1.65 4.785 1.255 4.905 1.255 4.905 1.315 4.845 1.315 4.845 1.65 5.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5.16 0.06 5.16 0.47 5.1 0.47 5.1 0.06 4.52 0.06 4.52 0.325 4.4 0.325 4.4 0.265 4.46 0.265 4.46 0.06 3.8 0.06 3.8 0.43 3.74 0.43 3.74 0.06 2.57 0.06 2.57 0.49 2.51 0.49 2.51 0.06 1.665 0.06 1.665 0.2 1.605 0.2 1.605 0.06 0.44 0.06 0.44 0.365 0.5 0.365 0.5 0.425 0.38 0.425 0.38 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.365 1.075 5.305 1.075 5.305 0.63 4.94 0.63 4.94 0.275 4.68 0.275 4.68 0.485 4.24 0.485 4.24 0.275 3.98 0.275 3.98 0.995 3.26 0.995 3.26 0.88 2.995 0.88 2.995 0.64 3.055 0.64 3.055 0.82 3.26 0.82 3.26 0.76 3.32 0.76 3.32 0.935 3.92 0.935 3.92 0.215 4.3 0.215 4.3 0.425 4.62 0.425 4.62 0.215 5 0.215 5 0.57 5.305 0.57 5.305 0.375 5.365 0.375 ;
      POLYGON 4.36 1.155 3.1 1.155 3.1 1.035 3.16 1.035 3.16 1.095 4.3 1.095 4.3 0.745 4.36 0.745 ;
      POLYGON 3.82 0.835 3.42 0.835 3.42 0.54 3.025 0.54 3.025 0.395 3.085 0.395 3.085 0.48 3.48 0.48 3.48 0.775 3.76 0.775 3.76 0.715 3.82 0.715 ;
      POLYGON 3.64 0.675 3.58 0.675 3.58 0.295 2.895 0.295 2.895 0.65 2.345 0.65 2.345 0.885 2.25 0.885 2.25 1.295 1.905 1.295 1.905 1.235 2.19 1.235 2.19 0.825 2.285 0.825 2.285 0.46 2.02 0.46 2.02 0.4 2.345 0.4 2.345 0.59 2.835 0.59 2.835 0.235 3.64 0.235 ;
      POLYGON 2.735 1.36 2.41 1.36 2.41 1.455 1.745 1.455 1.745 1.36 1.05 1.36 1.05 1.42 0.99 1.42 0.99 0.36 1.05 0.36 1.05 1.3 1.805 1.3 1.805 1.395 2.35 1.395 2.35 1.3 2.675 1.3 2.675 0.775 2.735 0.775 ;
      POLYGON 2.185 0.725 2.125 0.725 2.125 0.62 1.92 0.62 1.92 1.045 1.86 1.045 1.86 0.62 1.31 0.62 1.31 0.56 2.185 0.56 ;
      POLYGON 1.92 0.36 1.21 0.36 1.21 1.045 1.15 1.045 1.15 0.26 0.685 0.26 0.685 0.585 0.16 0.585 0.16 1.02 0.265 1.02 0.265 1.33 0.205 1.33 0.205 1.08 0.1 1.08 0.1 0.525 0.205 0.525 0.205 0.36 0.265 0.36 0.265 0.525 0.625 0.525 0.625 0.185 0.745 0.185 0.745 0.2 1.21 0.2 1.21 0.3 1.86 0.3 1.86 0.21 1.92 0.21 ;
  END
END MXI4X4

MACRO MXI4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MXI4XL 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9644 LAYER Metal1 ;
    ANTENNADIFFAREA 2.383925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0972 LAYER Metal1 ;
      ANTENNAMAXAREACAR 20.2098765 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 154.18209875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.215 1.02 0.135 1.02 0.135 0.73 0.06 0.73 0.06 0.6 0.135 0.6 0.135 0.54 0.215 0.54 ;
    END
  END Y
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.068 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.399177 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 15.0617285 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.435 0.815 3.935 0.895 ;
    END
  END S0
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.89 1.12 3.485 1.12 3.485 1.085 3.435 1.085 3.435 0.995 3.89 0.995 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.015 1.085 2.775 1.085 2.775 0.745 2.855 0.745 2.855 1.005 3.015 1.005 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.675 0.96 2.565 0.96 2.565 1.085 2.3 1.085 2.3 0.88 2.675 0.88 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.82 0.985 1.685 0.985 1.685 0.705 1.6 0.705 1.6 0.625 1.765 0.625 1.765 0.905 1.82 0.905 ;
    END
  END D
  PIN S1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 19.9074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.39 0.96 1.33 0.96 1.33 0.33 0.54 0.33 0.54 0.71 0.545 0.71 0.545 0.83 0.48 0.83 0.48 0.54 0.46 0.54 0.46 0.41 0.48 0.41 0.48 0.27 1.06 0.27 1.06 0.245 1.18 0.245 1.18 0.27 1.39 0.27 ;
    END
  END S1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 1.77 0 1.77 0 1.65 0.38 1.65 0.38 1.315 0.5 1.315 0.5 1.375 0.44 1.375 0.44 1.65 0.725 1.65 0.725 1.31 0.665 1.31 0.665 1.25 0.785 1.25 0.785 1.65 1.66 1.65 1.66 1.51 1.72 1.51 1.72 1.65 2.605 1.65 2.605 1.405 2.545 1.405 2.545 1.345 2.665 1.345 2.665 1.65 3.635 1.65 3.635 1.22 3.695 1.22 3.695 1.65 4.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 0.06 3.8 0.06 3.8 0.2 3.74 0.2 3.74 0.06 2.74 0.06 2.74 0.2 2.68 0.2 2.68 0.06 1.655 0.06 1.655 0.465 1.595 0.465 1.595 0.06 0.96 0.06 0.96 0.17 0.84 0.17 0.84 0.06 0.5 0.06 0.5 0.17 0.38 0.17 0.38 0.06 0 0.06 0 -0.06 4.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.095 1.185 4.05 1.185 4.05 1.245 3.99 1.245 3.99 1.125 4.035 1.125 4.035 0.36 3.58 0.36 3.58 0.24 3.175 0.24 3.175 1.04 3.115 1.04 3.115 0.36 2.52 0.36 2.52 0.22 2.04 0.22 2.04 0.855 1.92 0.855 1.92 0.795 1.98 0.795 1.98 0.16 2.58 0.16 2.58 0.3 3.115 0.3 3.115 0.18 3.64 0.18 3.64 0.3 4.095 0.3 ;
      POLYGON 3.335 1.305 3.275 1.305 3.275 1.245 2.36 1.245 2.36 1.37 1.82 1.37 1.82 1.35 1.55 1.35 1.55 1.41 1.49 1.41 1.49 1.29 1.88 1.29 1.88 1.31 2.3 1.31 2.3 1.185 3.275 1.185 3.275 0.395 3.335 0.395 ;
      POLYGON 3.015 0.645 2.38 0.645 2.38 0.78 2.3 0.78 2.3 0.565 3.015 0.565 ;
      POLYGON 2.36 0.46 2.2 0.46 2.2 1.15 2.075 1.15 2.075 1.21 2.015 1.21 2.015 1.15 1.39 1.15 1.39 1.38 0.885 1.38 0.885 1.32 1.33 1.32 1.33 1.09 2.14 1.09 2.14 0.4 2.36 0.4 ;
      POLYGON 1.23 1.21 1.17 1.21 1.17 1.15 0.315 1.15 0.315 0.74 0.375 0.74 0.375 1.09 1.17 1.09 1.17 0.63 1.11 0.63 1.11 0.57 1.23 0.57 ;
      POLYGON 1.07 0.985 0.76 0.985 0.76 0.99 0.585 0.99 0.585 0.93 0.7 0.93 0.7 0.63 0.64 0.63 0.64 0.57 0.76 0.57 0.76 0.925 1.01 0.925 1.01 0.865 1.07 0.865 ;
  END
END MXI4XL

MACRO NAND2BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX1 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.354275 LAYER Metal1 ;
    ANTENNADIFFAREA 0.5085 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.11196575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 102.15384625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.32 1.315 0.26 1.315 0.26 1.015 0.22 1.015 0.22 0.935 0.26 0.935 0.26 0.56 0.125 0.56 0.125 0.38 0.185 0.38 0.185 0.5 0.32 0.5 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.29629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.575 0.83 0.76 0.985 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.17948725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.055 0.62 0.15 0.835 ;
    END
  END B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 0.06 0.5 0.06 0.5 0.625 0.435 0.625 0.435 0.06 0 0.06 0 -0.06 0.8 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.77 0 1.77 0 1.65 0.065 1.65 0.065 1.51 0.185 1.51 0.185 1.65 0.465 1.65 0.465 1.195 0.525 1.195 0.525 1.65 0.8 1.65 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 0.73 0.745 0.46 0.745 0.46 1.055 0.73 1.055 0.73 1.315 0.67 1.315 0.67 1.12 0.4 1.12 0.4 0.685 0.67 0.685 0.67 0.52 0.73 0.52 ;
  END
END NAND2BX1

MACRO NAND2BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX2 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.77625 LAYER Metal1 ;
    ANTENNADIFFAREA 0.8432 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.26923075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 105.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.75 1.48 0.69 1.48 0.69 1.17 0.34 1.17 0.34 1.48 0.28 1.48 0.28 1.1 0.69 1.1 0.69 0.85 0.075 0.85 0.075 0.55 0.585 0.55 0.585 0.25 0.645 0.25 0.645 0.61 0.155 0.61 0.155 0.79 0.75 0.79 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.83333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 0.775 1.19 0.935 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 1.035 0.075 1.035 0.075 0.955 0.405 0.955 0.405 0.92 0.54 0.92 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.075 1.65 0.075 1.105 0.135 1.105 0.135 1.65 0.485 1.65 0.485 1.23 0.545 1.23 0.545 1.65 0.895 1.65 0.895 1.235 0.955 1.235 0.955 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 0.955 0.06 0.955 0.49 0.895 0.49 0.895 0.06 0.335 0.06 0.335 0.49 0.275 0.49 0.275 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.19 0.61 0.96 0.61 0.96 1.105 1.19 1.105 1.19 1.225 1.13 1.225 1.13 1.17 0.9 1.17 0.9 0.73 0.32 0.73 0.32 0.67 0.9 0.67 0.9 0.55 1.13 0.55 1.13 0.39 1.19 0.39 ;
  END
END NAND2BX2

MACRO NAND2BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BX4 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.30495 LAYER Metal1 ;
    ANTENNADIFFAREA 1.438 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.15341875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 89.69230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.565 1.48 1.505 1.48 1.505 1.15 1.155 1.15 1.155 1.48 1.095 1.48 1.095 1.15 0.745 1.15 0.745 1.48 0.685 1.48 0.685 1.15 0.335 1.15 0.335 1.48 0.275 1.48 0.275 1.09 1.445 1.09 1.445 0.86 0.065 0.86 0.065 0.545 0.145 0.545 0.145 0.55 0.685 0.55 0.685 0.25 0.745 0.25 0.745 0.55 1.305 0.55 1.305 0.25 1.365 0.25 1.365 0.61 0.145 0.61 0.145 0.8 1.505 0.8 1.505 1.09 1.565 1.09 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.602564 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.385 0.925 1.32 1.005 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.73 0.74 1.975 0.885 ;
    END
  END AN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.23 0.13 1.23 0.13 1.65 0.48 1.65 0.48 1.23 0.54 1.23 0.54 1.65 0.89 1.65 0.89 1.23 0.95 1.23 0.95 1.65 1.3 1.65 1.3 1.23 1.36 1.23 1.36 1.65 1.71 1.65 1.71 1.23 1.77 1.23 1.77 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 1.675 0.06 1.675 0.51 1.615 0.51 1.615 0.06 1.055 0.06 1.055 0.49 0.995 0.49 0.995 0.06 0.435 0.06 0.435 0.49 0.375 0.49 0.375 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.975 1.48 1.915 1.48 1.915 1.09 1.67 1.09 1.67 1.01 1.61 1.01 1.61 0.73 0.39 0.73 0.39 0.67 1.495 0.67 1.495 0.6 1.82 0.6 1.82 0.25 1.88 0.25 1.88 0.66 1.67 0.66 1.67 0.95 1.73 0.95 1.73 1.03 1.975 1.03 ;
  END
END NAND2BX4

MACRO NAND2BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2BXL 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.332 LAYER Metal1 ;
    ANTENNADIFFAREA 0.454525 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 20.49382725 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 172.31481475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.32 1.22 0.26 1.22 0.26 1.145 0.14 1.145 0.14 1.3 0.055 1.3 0.055 0.59 0.1 0.59 0.1 0.54 0.16 0.54 0.16 0.73 0.115 0.73 0.115 1.085 0.32 1.085 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.12962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 1.12 0.66 1.12 0.66 1.015 0.575 1.015 0.575 0.9 0.74 0.9 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.83333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.365 0.73 0.28 0.73 0.28 1.005 0.185 1.005 0.185 0.885 0.22 0.885 0.22 0.6 0.365 0.6 ;
    END
  END B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 0.06 0.525 0.06 0.525 0.635 0.465 0.635 0.465 0.06 0 0.06 0 -0.06 0.8 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.77 0 1.77 0 1.65 0.09 1.65 0.09 1.51 0.15 1.51 0.15 1.65 0.465 1.65 0.465 1.51 0.525 1.51 0.525 1.65 0.8 1.65 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 0.73 0.84 0.5 0.84 0.5 1.18 0.73 1.18 0.73 1.3 0.67 1.3 0.67 1.24 0.44 1.24 0.44 1.015 0.355 1.015 0.355 0.955 0.44 0.955 0.44 0.74 0.67 0.74 0.67 0.52 0.73 0.52 ;
  END
END NAND2BXL

MACRO NAND2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X1 0 0 ;
  SIZE 0.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2241 LAYER Metal1 ;
    ANTENNADIFFAREA 0.4392 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.555 0.9 0.335 0.9 0.335 1.34 0.275 1.34 0.275 0.84 0.435 0.84 0.435 0.315 0.495 0.315 0.495 0.76 0.555 0.76 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.025641 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.095 0.775 0.215 0.95 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.295 0.44 0.375 0.745 ;
    END
  END B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 0.06 0.13 0.06 0.13 0.555 0.07 0.555 0.07 0.06 0 0.06 0 -0.06 0.6 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.09 0.13 1.09 0.13 1.65 0.43 1.65 0.43 1.51 0.55 1.51 0.55 1.65 0.6 1.65 ;
    END
  END VDD
END NAND2X1

MACRO NAND2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X2 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4415 LAYER Metal1 ;
    ANTENNADIFFAREA 0.7417 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.95 0.995 0.745 0.995 0.745 1.34 0.685 1.34 0.685 0.99 0.335 0.99 0.335 1.34 0.275 1.34 0.275 0.93 0.89 0.93 0.89 0.84 0.87 0.84 0.87 0.76 0.89 0.76 0.89 0.56 0.455 0.56 0.455 0.315 0.515 0.315 0.515 0.495 0.95 0.495 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.69230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.37 0.64 0.62 0.72 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.5384615 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.81 0.86 0.07 0.86 0.07 0.78 0.22 0.78 0.22 0.675 0.28 0.675 0.28 0.78 0.75 0.78 0.75 0.625 0.81 0.625 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.885 0.06 0.885 0.435 0.765 0.435 0.765 0.06 0.205 0.06 0.205 0.565 0.145 0.565 0.145 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.98 0.13 0.98 0.13 1.65 0.45 1.65 0.45 1.085 0.57 1.085 0.57 1.65 0.83 1.65 0.83 1.51 0.96 1.51 0.96 1.65 1 1.65 ;
    END
  END VDD
END NAND2X2

MACRO NAND2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X4 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7344 LAYER Metal1 ;
    ANTENNADIFFAREA 1.3088 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.695 0.895 1.565 0.895 1.565 1.345 1.505 1.345 1.505 0.995 1.155 0.995 1.155 1.345 1.095 1.345 1.095 0.995 0.745 0.995 0.745 1.345 0.685 1.345 0.685 1 0.335 1 0.335 1.345 0.275 1.345 0.275 0.935 1.505 0.935 1.505 0.815 1.62 0.815 1.62 0.595 0.595 0.595 0.595 0.305 0.655 0.305 0.655 0.53 1.215 0.53 1.215 0.305 1.275 0.305 1.275 0.53 1.695 0.53 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.87179475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.23 0.875 0.58 0.875 0.58 0.815 0.995 0.815 0.995 0.795 1.075 0.795 1.075 0.815 1.23 0.815 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.74358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 0.715 0.17 0.715 0.17 0.625 0.3 0.625 0.3 0.655 1.54 0.655 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.615 0.06 1.615 0.43 1.555 0.43 1.555 0.06 0.965 0.06 0.965 0.43 0.905 0.43 0.905 0.06 0.345 0.06 0.345 0.545 0.285 0.545 0.285 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.955 0.13 0.955 0.13 1.65 0.48 1.65 0.48 1.105 0.54 1.105 0.54 1.65 0.89 1.65 0.89 1.105 0.95 1.105 0.95 1.65 1.3 1.65 1.3 1.105 1.36 1.105 1.36 1.65 1.71 1.65 1.71 0.965 1.77 0.965 1.77 1.65 2 1.65 ;
    END
  END VDD
END NAND2X4

MACRO NAND2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X6 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0308 LAYER Metal1 ;
    ANTENNADIFFAREA 1.9932 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.61 1.045 2.395 1.045 2.395 1.345 2.335 1.345 2.335 1.045 1.985 1.045 1.985 1.345 1.925 1.345 1.925 1.045 1.575 1.045 1.575 1.345 1.515 1.345 1.515 1.045 1.165 1.045 1.165 1.345 1.105 1.345 1.105 1.045 0.745 1.045 0.745 1.345 0.685 1.345 0.685 1.045 0.335 1.045 0.335 1.345 0.275 1.345 0.275 0.985 2.53 0.985 2.53 0.555 0.51 0.555 0.51 0.305 0.57 0.305 0.57 0.495 1.41 0.495 1.41 0.305 1.47 0.305 1.47 0.495 2.09 0.495 2.09 0.305 2.15 0.305 2.15 0.495 2.595 0.495 2.595 0.965 2.61 0.965 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.17505 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.97343625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.125 0.875 2.01 0.875 2.01 0.895 1.93 0.895 1.93 0.875 0.47 0.875 0.47 0.815 2.125 0.815 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.17505 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.361611 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.47 0.88 2.41 0.88 2.41 0.745 0.205 0.745 0.205 0.685 0.33 0.685 0.33 0.6 0.41 0.6 0.41 0.685 2.47 0.685 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 0.06 1.84 0.06 1.84 0.43 1.72 0.43 1.72 0.06 0.965 0.06 0.965 0.43 0.845 0.43 0.845 0.06 0.23 0.06 0.23 0.595 0.17 0.595 0.17 0.06 0 0.06 0 -0.06 2.8 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.955 0.13 0.955 0.13 1.65 0.48 1.65 0.48 1.105 0.54 1.105 0.54 1.65 0.9 1.65 0.9 1.105 0.96 1.105 0.96 1.65 1.31 1.65 1.31 1.105 1.37 1.105 1.37 1.65 1.72 1.65 1.72 1.105 1.78 1.105 1.78 1.65 2.13 1.65 2.13 1.105 2.19 1.105 2.19 1.65 2.54 1.65 2.54 1.105 2.6 1.105 2.6 1.65 2.8 1.65 ;
    END
  END VDD
END NAND2X6

MACRO NAND2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X8 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.203 LAYER Metal1 ;
    ANTENNADIFFAREA 2.4788 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.005 1.085 2.795 1.085 2.795 1.44 2.735 1.44 2.735 1.075 2.385 1.075 2.385 1.44 2.325 1.44 2.325 1.075 1.975 1.075 1.975 1.44 1.915 1.44 1.915 1.075 1.565 1.075 1.565 1.44 1.505 1.44 1.505 1.075 1.155 1.075 1.155 1.44 1.095 1.44 1.095 1.075 0.745 1.075 0.745 1.44 0.685 1.44 0.685 1.075 0.335 1.075 0.335 1.44 0.275 1.44 0.275 0.995 0.335 0.995 0.335 1.015 2.925 1.015 2.925 0.665 0.48 0.665 0.48 0.365 0.54 0.365 0.54 0.605 1.3 0.605 1.3 0.365 1.36 0.365 1.36 0.605 2.12 0.605 2.12 0.365 2.18 0.365 2.18 0.605 2.84 0.605 2.84 0.365 2.9 0.365 2.9 0.605 3.005 0.605 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.24967825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.865 0.925 0.45 0.925 0.45 0.865 2.615 0.865 2.615 0.815 2.72 0.815 2.72 0.865 2.865 0.865 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.19176325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.56 0.79 0.215 0.79 0.215 0.655 0.345 0.655 0.345 0.73 2.56 0.73 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 0.06 2.59 0.06 2.59 0.545 2.47 0.545 2.47 0.06 1.8 0.06 1.8 0.545 1.68 0.545 1.68 0.06 0.935 0.06 0.935 0.545 0.815 0.545 0.815 0.06 0.23 0.06 0.23 0.595 0.17 0.595 0.17 0.06 0 0.06 0 -0.06 3.2 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.995 0.13 0.995 0.13 1.65 0.48 1.65 0.48 1.2 0.54 1.2 0.54 1.65 0.89 1.65 0.89 1.2 0.95 1.2 0.95 1.65 1.3 1.65 1.3 1.2 1.36 1.2 1.36 1.65 1.71 1.65 1.71 1.2 1.77 1.2 1.77 1.65 2.12 1.65 2.12 1.2 2.18 1.2 2.18 1.65 2.53 1.65 2.53 1.2 2.59 1.2 2.59 1.65 2.94 1.65 2.94 1.2 3 1.2 3 1.65 3.2 1.65 ;
    END
  END VDD
END NAND2X8

MACRO NAND2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2XL 0 0 ;
  SIZE 0.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2052 LAYER Metal1 ;
    ANTENNADIFFAREA 0.34005 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 0.565 0.52 0.565 0.52 1.16 0.24 1.16 0.24 1.1 0.46 1.1 0.46 0.565 0.415 0.565 0.415 0.41 0.54 0.41 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.83333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.24 0.735 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.4 0.905 0.23 0.905 0.23 0.815 0.335 0.815 0.335 0.72 0.4 0.72 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.38 0.13 1.38 0.13 1.65 0.47 1.65 0.47 1.38 0.53 1.38 0.53 1.65 0.6 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 0.06 0.165 0.06 0.165 0.54 0.105 0.54 0.105 0.06 0 0.06 0 -0.06 0.6 -0.06 ;
    END
  END VSS
END NAND2XL

MACRO NAND3BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.574475 LAYER Metal1 ;
    ANTENNADIFFAREA 0.721475 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.640171 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 152.30769225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.615 1.48 0.555 1.48 0.555 1.14 0.205 1.14 0.205 1.48 0.145 1.48 0.145 1.2 0.085 1.2 0.085 1.12 0.115 1.12 0.115 0.485 0.2 0.485 0.2 0.32 0.26 0.32 0.26 0.56 0.18 0.56 0.18 1.08 0.615 1.08 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.12962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.78 0.94 1.085 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.923077 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.62 0.54 1.02 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.923077 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.62 0.34 1.02 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.35 1.65 0.35 1.2 0.41 1.2 0.41 1.65 0.76 1.65 0.76 1.2 0.82 1.2 0.82 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.775 0.06 0.775 0.56 0.715 0.56 0.715 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.06 1.21 1 1.21 1 0.7 0.73 0.7 0.73 0.835 0.67 0.835 0.67 0.64 0.95 0.64 0.95 0.46 1.01 0.46 1.01 0.64 1.06 0.64 ;
  END
END NAND3BX1

MACRO NAND3BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.908 LAYER Metal1 ;
    ANTENNADIFFAREA 1.22005 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 15.5213675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 120.102564 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.26 1.345 1.2 1.345 1.2 1.125 0.85 1.125 0.85 1.345 0.79 1.345 0.79 1.125 0.43 1.125 0.43 1.345 0.37 1.345 0.37 1.085 0.15 1.085 0.15 0.335 0.825 0.335 0.825 0.395 0.21 0.395 0.21 1.005 0.43 1.005 0.43 1.065 1.2 1.065 1.2 1.02 1.26 1.02 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.96 0.965 0.88 0.965 0.88 0.895 0.53 0.895 0.53 0.815 0.96 0.815 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.79487175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 0.92 1.06 0.92 1.06 0.715 0.47 0.715 0.47 0.655 1.13 0.655 1.13 0.715 1.14 0.715 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.57 0.92 1.54 0.92 1.54 1.125 1.46 1.125 1.46 0.785 1.49 0.785 1.49 0.655 1.57 0.655 ;
    END
  END AN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.165 1.65 0.165 1.225 0.225 1.225 0.225 1.65 0.575 1.65 0.575 1.225 0.635 1.225 0.635 1.65 0.995 1.65 0.995 1.225 1.055 1.225 1.055 1.65 1.405 1.65 1.405 1.225 1.465 1.225 1.465 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.38 0.06 1.38 0.335 1.44 0.335 1.44 0.395 1.32 0.395 1.32 0.06 0.295 0.06 0.295 0.17 0.175 0.17 0.175 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.73 1.075 1.67 1.075 1.67 0.555 1.335 0.555 1.335 0.76 1.275 0.76 1.275 0.555 0.37 0.555 0.37 0.735 0.31 0.735 0.31 0.495 1.585 0.495 1.585 0.435 1.645 0.435 1.645 0.495 1.73 0.495 ;
  END
END NAND3BX2

MACRO NAND3BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BX4 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5701 LAYER Metal1 ;
    ANTENNADIFFAREA 2.1865 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.419658 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 103.64102575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.41 1.425 2.35 1.425 2.35 1.185 2 1.185 2 1.425 1.94 1.425 1.94 1.185 1.59 1.185 1.59 1.425 1.53 1.425 1.53 1.185 1.18 1.185 1.18 1.425 1.12 1.425 1.12 1.185 0.77 1.185 0.77 1.425 0.71 1.425 0.71 1.185 0.36 1.185 0.36 1.425 0.3 1.425 0.3 1.095 0.08 1.095 0.08 0.54 0.06 0.54 0.06 0.41 1.95 0.41 1.95 0.47 0.14 0.47 0.14 1.035 0.36 1.035 0.36 1.125 2.41 1.125 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.70512825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.265 0.865 1.605 0.865 1.605 0.805 1.285 0.805 1.285 0.865 0.66 0.865 0.66 0.715 0.4 0.715 0.4 0.655 0.435 0.655 0.435 0.625 0.565 0.625 0.565 0.655 0.72 0.655 0.72 0.805 1.225 0.805 1.225 0.745 1.665 0.745 1.665 0.805 2.265 0.805 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.775 0.795 2.485 0.795 2.485 0.705 2.365 0.705 2.365 0.625 2.565 0.625 2.565 0.715 2.775 0.715 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.24358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.885 0.705 1.765 0.705 1.765 0.645 1.125 0.645 1.125 0.705 0.82 0.705 0.82 0.645 0.835 0.645 0.835 0.625 0.965 0.625 0.965 0.645 1.065 0.645 1.065 0.585 1.825 0.585 1.825 0.645 1.885 0.645 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.77 0 1.77 0 1.65 0.095 1.65 0.095 1.305 0.155 1.305 0.155 1.65 0.505 1.65 0.505 1.305 0.565 1.305 0.565 1.65 0.915 1.65 0.915 1.305 0.975 1.305 0.975 1.65 1.325 1.65 1.325 1.305 1.385 1.305 1.385 1.65 1.735 1.65 1.735 1.305 1.795 1.305 1.795 1.65 2.145 1.65 2.145 1.305 2.205 1.305 2.205 1.65 2.555 1.65 2.555 1.055 2.615 1.055 2.615 1.65 3 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 0.06 2.56 0.06 2.56 0.435 2.5 0.435 2.5 0.06 1.315 0.06 1.315 0.16 1.375 0.16 1.375 0.22 1.255 0.22 1.255 0.06 0.165 0.06 0.165 0.16 0.225 0.16 0.225 0.22 0.105 0.22 0.105 0.06 0 0.06 0 -0.06 3 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.935 0.955 2.85 0.955 2.85 1.425 2.76 1.425 2.76 0.955 2.455 0.955 2.455 1.025 0.5 1.025 0.5 0.935 0.24 0.935 0.24 0.815 0.3 0.815 0.3 0.875 0.56 0.875 0.56 0.965 1.385 0.965 1.385 0.905 1.505 0.905 1.505 0.965 2.395 0.965 2.395 0.895 2.875 0.895 2.875 0.575 2.705 0.575 2.705 0.455 2.765 0.455 2.765 0.515 2.935 0.515 ;
  END
END NAND3BX4

MACRO NAND3BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3BXL 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4557 LAYER Metal1 ;
    ANTENNADIFFAREA 0.5536 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 28.12962975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 206.4814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 1.18 0.14 1.18 0.14 1.305 0.06 1.305 0.06 0.495 0.085 0.495 0.085 0.435 0.145 0.435 0.145 0.555 0.12 0.555 0.12 1.09 0.13 1.09 0.13 1.12 0.56 1.12 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.611111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.635 0.8 0.79 1.11 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.375 0.79 0.54 0.985 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.9444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.365 0.73 0.27 0.73 0.27 0.79 0.18 0.79 0.18 0.615 0.235 0.615 0.235 0.6 0.365 0.6 ;
    END
  END C
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.72 0.06 0.72 0.555 0.66 0.555 0.66 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.49 0.4 1.49 0.4 1.65 0.605 1.65 0.605 1.49 0.725 1.49 0.725 1.65 1 1.65 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 0.93 1.21 0.87 1.21 0.87 0.72 0.555 0.72 0.555 0.66 0.865 0.66 0.865 0.46 0.925 0.46 0.925 0.66 0.93 0.66 ;
  END
END NAND3BXL

MACRO NAND3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X1 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3252 LAYER Metal1 ;
    ANTENNADIFFAREA 0.6209 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.765 1.49 0.685 1.49 0.685 1.3 0.635 1.3 0.635 1.175 0.335 1.175 0.335 1.48 0.275 1.48 0.275 1.115 0.685 1.115 0.685 0.65 0.65 0.65 0.65 0.38 0.685 0.38 0.685 0.375 0.745 0.375 0.745 1.16 0.765 1.16 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.69230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.59 0.8 0.5 0.8 0.5 0.73 0.435 0.73 0.435 0.595 0.59 0.595 ;
    END
  END C
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.3846155 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.92 0.19 1.12 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.12820525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.41 0.945 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.2 0.13 1.2 0.13 1.65 0.48 1.65 0.48 1.24 0.54 1.24 0.54 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.13 0.06 0.13 0.62 0.07 0.62 0.07 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NAND3X1

MACRO NAND3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X2 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5415 LAYER Metal1 ;
    ANTENNADIFFAREA 1.0842 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.565 1.115 1.25 1.115 1.25 1.335 1.19 1.335 1.19 1.115 0.84 1.115 0.84 1.335 0.78 1.335 0.78 1.115 0.43 1.115 0.43 1.335 0.36 1.335 0.36 1.055 1.435 1.055 1.435 1.005 1.505 1.005 1.505 0.395 0.795 0.395 0.795 0.335 1.565 0.335 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.96 0.895 0.765 0.895 0.765 0.955 0.52 0.955 0.52 0.815 0.96 0.815 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.79487175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 0.92 1.06 0.92 1.06 0.715 0.47 0.715 0.47 0.655 1.14 0.655 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.3 0.735 1.24 0.735 1.24 0.555 0.37 0.555 0.37 0.735 0.26 0.735 0.26 0.6 0.31 0.6 0.31 0.495 1.3 0.495 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.165 1.65 0.165 0.945 0.225 0.945 0.225 1.65 0.575 1.65 0.575 1.215 0.635 1.215 0.635 1.65 0.985 1.65 0.985 1.215 1.045 1.215 1.045 1.65 1.395 1.65 1.395 1.215 1.455 1.215 1.455 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.435 0.06 1.435 0.17 1.315 0.17 1.315 0.06 0.265 0.06 0.265 0.335 0.325 0.335 0.325 0.395 0.205 0.395 0.205 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NAND3X2

MACRO NAND3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X4 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8904 LAYER Metal1 ;
    ANTENNADIFFAREA 2.015 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.74 1.11 2.525 1.11 2.525 1.405 2.465 1.405 2.465 1.185 2.115 1.185 2.115 1.405 2.055 1.405 2.055 1.185 1.705 1.185 1.705 1.405 1.645 1.405 1.645 1.185 1.295 1.185 1.295 1.405 1.235 1.405 1.235 1.185 0.885 1.185 0.885 1.405 0.825 1.405 0.825 1.185 0.475 1.185 0.475 1.405 0.415 1.405 0.415 1.015 0.475 1.015 0.475 1.125 2.465 1.125 2.465 1.04 2.525 1.04 2.525 1.05 2.66 1.05 2.66 0.98 2.68 0.98 2.68 0.465 0.895 0.465 0.895 0.405 2.74 0.405 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.0641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.555 0.94 2.365 0.94 2.365 1.025 0.64 1.025 0.64 0.915 0.305 0.915 0.305 0.895 0.235 0.895 0.235 0.815 0.365 0.815 0.365 0.855 0.7 0.855 0.7 0.965 1.475 0.965 1.475 0.885 1.595 0.885 1.595 0.965 2.305 0.965 2.305 0.88 2.495 0.88 2.495 0.82 2.555 0.82 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.19230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.395 0.745 2.205 0.745 2.205 0.865 1.695 0.865 1.695 0.785 1.325 0.785 1.325 0.865 0.8 0.865 0.8 0.755 0.515 0.755 0.515 0.695 0.86 0.695 0.86 0.805 1.265 0.805 1.265 0.725 1.755 0.725 1.755 0.805 2.145 0.805 2.145 0.685 2.26 0.685 2.26 0.6 2.34 0.6 2.34 0.625 2.395 0.625 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.19230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.985 0.705 1.855 0.705 1.855 0.625 1.165 0.625 1.165 0.705 0.96 0.705 0.96 0.645 1.035 0.645 1.035 0.565 1.915 0.565 1.915 0.645 1.985 0.645 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 1.77 0 1.77 0 1.65 0.21 1.65 0.21 1.015 0.27 1.015 0.27 1.65 0.62 1.65 0.62 1.285 0.68 1.285 0.68 1.65 1.03 1.65 1.03 1.285 1.09 1.285 1.09 1.65 1.44 1.65 1.44 1.285 1.5 1.285 1.5 1.65 1.85 1.65 1.85 1.285 1.91 1.285 1.91 1.65 2.26 1.65 2.26 1.285 2.32 1.285 2.32 1.65 2.67 1.65 2.67 1.285 2.73 1.285 2.73 1.65 2.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 0.06 2.63 0.06 2.63 0.16 2.69 0.16 2.69 0.22 2.57 0.22 2.57 0.06 1.455 0.06 1.455 0.16 1.515 0.16 1.515 0.22 1.395 0.22 1.395 0.06 0.37 0.06 0.37 0.435 0.31 0.435 0.31 0.06 0 0.06 0 -0.06 2.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NAND3X4

MACRO NAND3X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X6 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.305 LAYER Metal1 ;
    ANTENNADIFFAREA 3.0999 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.14 1.24 3.895 1.24 3.895 1.43 3.835 1.43 3.835 1.24 3.485 1.24 3.485 1.3 3.425 1.3 3.425 1.24 3.075 1.24 3.075 1.3 3.015 1.3 3.015 1.24 2.665 1.24 2.665 1.43 2.605 1.43 2.605 1.24 2.23 1.24 2.23 1.3 2.17 1.3 2.17 1.24 1.68 1.24 1.68 1.3 1.62 1.3 1.62 1.24 1.27 1.24 1.27 1.3 1.21 1.3 1.21 1.24 0.86 1.24 0.86 1.3 0.8 1.3 0.8 1.24 0.45 1.24 0.45 1.3 0.39 1.3 0.39 1.18 2.605 1.18 2.605 1.07 2.665 1.07 2.665 1.18 4.06 1.18 4.06 0.98 4.08 0.98 4.08 0.6 3.405 0.6 3.405 0.49 2.025 0.49 2.025 0.6 1.965 0.6 1.965 0.38 0.835 0.38 0.835 0.6 0.775 0.6 0.775 0.32 2.025 0.32 2.025 0.43 3.405 0.43 3.405 0.32 3.465 0.32 3.465 0.54 4.14 0.54 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.17505 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.866324 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.97 0.88 3.96 0.88 3.96 1.08 2.925 1.08 2.925 0.97 2.505 0.97 2.505 1.08 0.345 1.08 0.345 0.895 0.235 0.895 0.235 0.815 0.405 0.815 0.405 1.02 1.425 1.02 1.425 0.91 1.545 0.91 1.545 1.02 2.445 1.02 2.445 0.91 2.985 0.91 2.985 1.02 3.9 1.02 3.9 0.76 3.97 0.76 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.17505 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.61525275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.795 0.92 3.085 0.92 3.085 0.81 2.345 0.81 2.345 0.92 1.645 0.92 1.645 0.81 1.325 0.81 1.325 0.865 1.165 0.865 1.165 0.92 0.505 0.92 0.505 0.86 1.105 0.86 1.105 0.805 1.265 0.805 1.265 0.75 1.705 0.75 1.705 0.86 2.285 0.86 2.285 0.75 3.145 0.75 3.145 0.86 3.66 0.86 3.66 0.79 3.74 0.79 3.74 0.86 3.795 0.86 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.17505 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.192802 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.415 0.76 3.245 0.76 3.245 0.65 2.185 0.65 2.185 0.76 1.805 0.76 1.805 0.65 1.165 0.65 1.165 0.705 1.005 0.705 1.005 0.76 0.885 0.76 0.885 0.7 0.945 0.7 0.945 0.625 1.105 0.625 1.105 0.59 1.865 0.59 1.865 0.7 2.125 0.7 2.125 0.59 3.305 0.59 3.305 0.7 3.415 0.7 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 1.77 0 1.77 0 1.65 0.185 1.65 0.185 1.04 0.245 1.04 0.245 1.65 0.565 1.65 0.565 1.34 0.685 1.34 0.685 1.4 0.625 1.4 0.625 1.65 0.975 1.65 0.975 1.34 1.095 1.34 1.095 1.4 1.035 1.4 1.035 1.65 1.385 1.65 1.385 1.34 1.505 1.34 1.505 1.4 1.445 1.4 1.445 1.65 1.795 1.65 1.795 1.34 1.915 1.34 1.915 1.4 1.855 1.4 1.855 1.65 2.345 1.65 2.345 1.34 2.465 1.34 2.465 1.4 2.405 1.4 2.405 1.65 2.78 1.65 2.78 1.34 2.9 1.34 2.9 1.4 2.84 1.4 2.84 1.65 3.19 1.65 3.19 1.34 3.31 1.34 3.31 1.4 3.25 1.4 3.25 1.65 3.6 1.65 3.6 1.34 3.72 1.34 3.72 1.4 3.66 1.4 3.66 1.65 4.01 1.65 4.01 1.34 4.13 1.34 4.13 1.4 4.07 1.4 4.07 1.65 4.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 0.06 2.81 0.06 2.81 0.16 2.87 0.16 2.87 0.22 2.75 0.22 2.75 0.06 1.43 0.06 1.43 0.16 1.49 0.16 1.49 0.22 1.37 0.22 1.37 0.06 0.345 0.06 0.345 0.63 0.285 0.63 0.285 0.06 0 0.06 0 -0.06 4.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NAND3X6

MACRO NAND3X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3X8 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.12375 LAYER Metal1 ;
    ANTENNADIFFAREA 3.849075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.625 1.46 4.525 1.46 4.525 1.11 4.175 1.11 4.175 1.46 4.115 1.46 4.115 1.27 3.765 1.27 3.765 1.46 3.705 1.46 3.705 1.27 3.32 1.27 3.32 1.33 3.26 1.33 3.26 1.27 2.91 1.27 2.91 1.33 2.85 1.33 2.85 1.27 2.5 1.27 2.5 1.33 2.44 1.33 2.44 1.27 2.085 1.27 2.085 1.33 2.025 1.33 2.025 1.27 1.64 1.27 1.64 1.46 1.58 1.46 1.58 1.27 1.23 1.27 1.23 1.33 1.17 1.33 1.17 1.27 0.82 1.27 0.82 1.33 0.76 1.33 0.76 1.27 0.375 1.27 0.375 1.46 0.315 1.46 0.315 1.195 0.375 1.195 0.375 1.21 1.58 1.21 1.58 1.06 1.64 1.06 1.64 1.21 3.705 1.21 3.705 1.06 3.765 1.06 3.765 1.21 4.115 1.21 4.115 1.015 4.175 1.015 4.175 1.05 4.46 1.05 4.46 0.98 4.565 0.98 4.565 0.465 0.775 0.465 0.775 0.405 4.625 0.405 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.952381 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.86 0.945 3.79 0.945 3.79 0.96 3.605 0.96 3.605 1.11 1.74 1.11 1.74 0.96 1.34 0.96 1.34 1.11 0.475 1.11 0.475 1.095 0.28 1.095 0.28 0.92 0.26 0.92 0.26 0.79 0.34 0.79 0.34 1.035 0.535 1.035 0.535 1.05 1.28 1.05 1.28 0.885 1.4 0.885 1.4 0.9 1.8 0.9 1.8 1.05 2.61 1.05 2.61 0.945 2.55 0.945 2.55 0.885 2.67 0.885 2.67 1.05 3.545 1.05 3.545 0.9 3.73 0.9 3.73 0.885 3.86 0.885 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.18404125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.245 0.895 4.035 0.895 4.035 0.785 3.63 0.785 3.63 0.8 3.445 0.8 3.445 0.95 2.97 0.95 2.97 0.8 2.77 0.8 2.77 0.785 2.4 0.785 2.4 0.8 2.34 0.8 2.34 0.95 1.9 0.95 1.9 0.8 1.5 0.8 1.5 0.785 1.1 0.785 1.1 0.95 0.635 0.95 0.635 0.935 0.45 0.935 0.45 0.875 0.695 0.875 0.695 0.89 1.04 0.89 1.04 0.725 1.56 0.725 1.56 0.74 1.96 0.74 1.96 0.89 2.28 0.89 2.28 0.74 2.34 0.74 2.34 0.725 2.83 0.725 2.83 0.74 3.03 0.74 3.03 0.89 3.385 0.89 3.385 0.74 3.51 0.74 3.51 0.725 4.245 0.725 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.81724575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.465 0.8 4.345 0.8 4.345 0.625 3.285 0.625 3.285 0.79 3.165 0.79 3.165 0.73 3.225 0.73 3.225 0.625 2.12 0.625 2.12 0.73 2.18 0.73 2.18 0.79 2.06 0.79 2.06 0.625 0.94 0.625 0.94 0.79 0.795 0.79 0.795 0.73 0.86 0.73 0.86 0.6 0.88 0.6 0.88 0.565 4.405 0.565 4.405 0.74 4.465 0.74 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.11 1.65 0.11 1.02 0.17 1.02 0.17 1.65 0.525 1.65 0.525 1.37 0.645 1.37 0.645 1.43 0.585 1.43 0.585 1.65 0.935 1.65 0.935 1.37 1.055 1.37 1.055 1.43 0.995 1.43 0.995 1.65 1.345 1.65 1.345 1.37 1.465 1.37 1.465 1.43 1.405 1.43 1.405 1.65 1.755 1.65 1.755 1.37 1.875 1.37 1.875 1.43 1.815 1.43 1.815 1.65 2.2 1.65 2.2 1.37 2.32 1.37 2.32 1.43 2.26 1.43 2.26 1.65 2.615 1.65 2.615 1.37 2.735 1.37 2.735 1.43 2.675 1.43 2.675 1.65 3.025 1.65 3.025 1.37 3.145 1.37 3.145 1.43 3.085 1.43 3.085 1.65 3.435 1.65 3.435 1.37 3.555 1.37 3.555 1.43 3.495 1.43 3.495 1.65 3.88 1.65 3.88 1.37 4 1.37 4 1.43 3.94 1.43 3.94 1.65 4.29 1.65 4.29 1.37 4.41 1.37 4.41 1.43 4.35 1.43 4.35 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 3.97 0.06 3.97 0.17 3.85 0.17 3.85 0.06 2.765 0.06 2.765 0.17 2.645 0.17 2.645 0.06 1.395 0.06 1.395 0.17 1.275 0.17 1.275 0.06 0.305 0.06 0.305 0.485 0.245 0.485 0.245 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NAND3X8

MACRO NAND3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3XL 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3156 LAYER Metal1 ;
    ANTENNADIFFAREA 0.4939 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 1.225 0.86 1.225 0.86 1.165 0.405 1.165 0.405 1.105 0.86 1.105 0.86 0.98 0.87 0.98 0.87 0.54 0.94 0.54 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.755 0.88 0.66 0.88 0.66 0.395 0.74 0.395 0.74 0.76 0.755 0.76 ;
    END
  END C
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.34 1.005 0.03 1.005 0.03 0.735 0.11 0.735 0.11 0.79 0.34 0.79 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 0.89 0.48 0.89 0.48 0.54 0.46 0.54 0.46 0.41 0.54 0.41 0.54 0.48 0.56 0.48 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.23 1.65 0.23 1.105 0.29 1.105 0.29 1.65 0.6 1.65 0.6 1.51 0.66 1.51 0.66 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.29 0.06 0.29 0.635 0.23 0.635 0.23 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NAND3XL

MACRO NAND4BBX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX1 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.958325 LAYER Metal1 ;
    ANTENNADIFFAREA 1.20715 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.381624 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 126.30769225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.345 1.085 1.34 1.085 1.34 1.48 1.28 1.48 1.28 1.26 0.91 1.26 0.91 1.48 0.85 1.48 0.85 1.2 1.26 1.2 1.26 0.98 1.285 0.98 1.285 0.365 0.615 0.365 0.615 0.305 1.345 0.305 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.735 0.705 0.565 0.705 0.565 0.905 0.435 0.905 0.435 0.815 0.485 0.815 0.485 0.625 0.735 0.625 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 1.1 0.835 1.1 0.835 0.625 0.915 0.625 0.915 0.79 0.94 0.79 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.765 1.225 1.685 1.225 1.685 0.895 1.635 0.895 1.635 0.815 1.675 0.815 1.675 0.775 1.765 0.775 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.175 1.035 0.06 1.035 0.06 0.73 0.03 0.73 0.03 0.6 0.14 0.6 0.14 0.88 0.175 0.88 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.135 0.13 1.135 0.13 1.65 0.645 1.65 0.645 1.36 0.705 1.36 0.705 1.65 1.055 1.65 1.055 1.36 1.115 1.36 1.115 1.65 1.485 1.65 1.485 1.09 1.545 1.09 1.545 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.505 0.06 1.505 0.395 1.445 0.395 1.445 0.06 0.13 0.06 0.13 0.5 0.07 0.5 0.07 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.925 1.21 1.865 1.21 1.865 0.675 1.575 0.675 1.575 0.69 1.455 0.69 1.455 0.63 1.515 0.63 1.515 0.615 1.75 0.615 1.75 0.415 1.81 0.415 1.81 0.615 1.925 0.615 ;
      POLYGON 1.185 0.665 1.04 0.665 1.04 0.525 0.335 0.525 0.335 1.16 0.275 1.16 0.275 0.405 0.335 0.405 0.335 0.465 1.1 0.465 1.1 0.605 1.185 0.605 ;
  END
END NAND4BBX1

MACRO NAND4BBX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX2 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.69135 LAYER Metal1 ;
    ANTENNADIFFAREA 1.914425 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.455983 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 113.64102575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.925 1.155 2.88 1.155 2.88 1.375 2.82 1.375 2.82 1.155 2.43 1.155 2.43 1.375 2.37 1.375 2.37 1.155 2.02 1.155 2.02 1.375 1.96 1.375 1.96 1.155 1.61 1.155 1.61 1.375 1.55 1.375 1.55 1.005 1.765 1.005 1.765 1.095 2.865 1.095 2.865 0.44 2.925 0.44 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.765 0.995 2.685 0.995 2.685 0.73 2.66 0.73 2.66 0.52 2.74 0.52 2.74 0.65 2.765 0.65 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.54 0.995 2.25 0.995 2.25 0.705 2.33 0.705 2.33 0.79 2.54 0.79 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.795 1.165 0.565 1.165 0.565 0.815 0.65 0.815 0.65 1.005 0.795 1.005 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.465 1.165 0.385 1.165 0.385 0.895 0.235 0.895 0.235 0.815 0.465 0.815 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 1.77 0 1.77 0 1.65 0.46 1.65 0.46 1.265 0.52 1.265 0.52 1.65 1.345 1.65 1.345 1.005 1.405 1.005 1.405 1.65 1.755 1.65 1.755 1.255 1.815 1.255 1.815 1.65 2.165 1.65 2.165 1.255 2.225 1.255 2.225 1.65 2.575 1.65 2.575 1.255 2.635 1.255 2.635 1.65 3.025 1.65 3.025 0.985 3.085 0.985 3.085 1.65 3.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 0.06 1.51 0.06 1.51 0.415 1.39 0.415 1.39 0.355 1.45 0.355 1.45 0.06 0.545 0.06 0.545 0.555 0.485 0.555 0.485 0.06 0 0.06 0 -0.06 3.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.13 0.42 3.07 0.42 3.07 0.34 2.72 0.34 2.72 0.42 2.66 0.42 2.66 0.34 2.31 0.34 2.31 0.42 2.25 0.42 2.25 0.28 3.13 0.28 ;
      POLYGON 2.515 0.605 1.93 0.605 1.93 0.585 1.845 0.585 1.845 0.465 1.905 0.465 1.905 0.525 1.98 0.525 1.98 0.545 2.455 0.545 2.455 0.44 2.515 0.44 ;
      POLYGON 2.11 0.445 2.05 0.445 2.05 0.365 1.73 0.365 1.73 0.415 1.67 0.415 1.67 0.575 1.215 0.575 1.215 0.455 1.275 0.455 1.275 0.515 1.61 0.515 1.61 0.355 1.67 0.355 1.67 0.305 2.11 0.305 ;
      POLYGON 1.86 0.745 1.055 0.745 1.055 0.365 0.705 0.365 0.705 0.715 0.135 0.715 0.135 1.17 0.285 1.17 0.285 1.29 0.225 1.29 0.225 1.23 0.075 1.23 0.075 0.655 0.255 0.655 0.255 0.465 0.315 0.465 0.315 0.655 0.645 0.655 0.645 0.305 1.115 0.305 1.115 0.685 1.86 0.685 ;
      POLYGON 1.435 0.905 0.955 0.905 0.955 1.325 0.725 1.325 0.725 1.385 0.665 1.385 0.665 1.265 0.895 1.265 0.895 0.585 0.805 0.585 0.805 0.465 0.865 0.465 0.865 0.525 0.955 0.525 0.955 0.845 1.435 0.845 ;
  END
END NAND4BBX2

MACRO NAND4BBX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBX4 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.490975 LAYER Metal1 ;
    ANTENNADIFFAREA 3.2087 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.234 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.64519225 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 83.602564 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.325 0.56 3.915 0.56 3.915 1.085 4.195 1.085 4.195 1.365 4.135 1.365 4.135 1.145 3.785 1.145 3.785 1.365 3.725 1.365 3.725 1.145 3.375 1.145 3.375 1.365 3.315 1.365 3.315 1.145 2.965 1.145 2.965 1.365 2.905 1.365 2.905 1.145 2.555 1.145 2.555 1.365 2.495 1.365 2.495 1.145 2.145 1.145 2.145 1.365 2.085 1.365 2.085 1.145 1.735 1.145 1.735 1.365 1.675 1.365 1.675 1.145 1.325 1.145 1.325 1.365 1.265 1.365 1.265 1.005 1.565 1.005 1.565 1.085 3.855 1.085 3.855 0.42 3.915 0.42 3.915 0.5 4.265 0.5 4.265 0.42 4.325 0.42 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.755 0.985 3.675 0.985 3.675 0.73 3.66 0.73 3.66 0.5 3.74 0.5 3.74 0.65 3.755 0.65 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.14 0.985 2.84 0.985 2.84 0.705 2.92 0.705 2.92 0.74 3.14 0.74 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.76 0.54 1.26 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.76 0.34 1.26 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.77 0 1.77 0 1.65 0.405 1.65 0.405 1.36 0.465 1.36 0.465 1.65 1.06 1.65 1.06 1.005 1.12 1.005 1.12 1.65 1.47 1.65 1.47 1.245 1.53 1.245 1.53 1.65 1.88 1.65 1.88 1.245 1.94 1.245 1.94 1.65 2.29 1.65 2.29 1.245 2.35 1.245 2.35 1.65 2.7 1.65 2.7 1.245 2.76 1.245 2.76 1.65 3.11 1.65 3.11 1.245 3.17 1.245 3.17 1.65 3.52 1.65 3.52 1.245 3.58 1.245 3.58 1.65 3.93 1.65 3.93 1.245 3.99 1.245 3.99 1.65 4.34 1.65 4.34 0.975 4.4 0.975 4.4 1.65 4.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 0.06 1.68 0.06 1.68 0.415 1.56 0.415 1.56 0.355 1.62 0.355 1.62 0.06 1.21 0.06 1.21 0.355 1.27 0.355 1.27 0.415 1.15 0.415 1.15 0.06 0.39 0.06 0.39 0.5 0.33 0.5 0.33 0.06 0 0.06 0 -0.06 4.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.53 0.4 4.47 0.4 4.47 0.32 4.12 0.32 4.12 0.4 4.06 0.4 4.06 0.32 3.71 0.32 3.71 0.4 3.65 0.4 3.65 0.32 3.3 0.32 3.3 0.4 3.24 0.4 3.24 0.32 2.89 0.32 2.89 0.4 2.83 0.4 2.83 0.26 4.53 0.26 ;
      POLYGON 3.505 0.605 2.1 0.605 2.1 0.585 2.015 0.585 2.015 0.465 2.075 0.465 2.075 0.525 2.15 0.525 2.15 0.545 2.425 0.545 2.425 0.465 2.485 0.465 2.485 0.545 3.035 0.545 3.035 0.42 3.095 0.42 3.095 0.545 3.445 0.545 3.445 0.42 3.505 0.42 ;
      POLYGON 2.69 0.445 2.63 0.445 2.63 0.365 2.28 0.365 2.28 0.445 2.22 0.445 2.22 0.365 1.9 0.365 1.9 0.415 1.84 0.415 1.84 0.575 0.975 0.575 0.975 0.455 1.035 0.455 1.035 0.515 1.385 0.515 1.385 0.455 1.445 0.455 1.445 0.515 1.78 0.515 1.78 0.355 1.84 0.355 1.84 0.305 2.69 0.305 ;
      POLYGON 2.03 0.745 0.81 0.745 0.81 0.42 0.55 0.42 0.55 0.66 0.16 0.66 0.16 1.36 0.26 1.36 0.26 1.48 0.2 1.48 0.2 1.42 0.1 1.42 0.1 0.605 0.125 0.605 0.125 0.52 0.185 0.52 0.185 0.6 0.49 0.6 0.49 0.36 0.87 0.36 0.87 0.685 2.03 0.685 ;
      POLYGON 1.205 0.905 0.71 0.905 0.71 1.13 0.7 1.13 0.7 1.48 0.64 1.48 0.64 1.09 0.65 1.09 0.65 0.52 0.71 0.52 0.71 0.845 1.205 0.845 ;
  END
END NAND4BBX4

MACRO NAND4BBXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BBXL 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.88345 LAYER Metal1 ;
    ANTENNADIFFAREA 0.901675 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 27.26697525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 209.537037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.175 1.385 1.115 1.385 1.115 1.29 0.75 1.29 0.75 1.385 0.69 1.385 0.69 1.23 1.06 1.23 1.06 0.98 1.115 0.98 1.115 0.42 0.555 0.42 0.555 0.36 1.175 0.36 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.815 0.7 1.13 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 0.92 0.88 0.92 0.88 1.13 0.8 1.13 0.8 0.84 0.86 0.84 0.86 0.69 0.94 0.69 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.565 1.105 1.415 1.105 1.415 0.895 1.275 0.895 1.275 0.815 1.565 0.815 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.175 0.965 0.095 0.965 0.095 0.745 0.06 0.745 0.06 0.5 0.14 0.5 0.14 0.625 0.175 0.625 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.065 0.13 1.065 0.13 1.65 0.485 1.65 0.485 1.36 0.545 1.36 0.545 1.65 0.865 1.65 0.865 1.39 0.985 1.39 0.985 1.45 0.925 1.45 0.925 1.65 1.37 1.65 1.37 1.36 1.43 1.36 1.43 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.43 0.06 1.43 0.425 1.37 0.425 1.37 0.06 0.13 0.06 0.13 0.4 0.07 0.4 0.07 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.725 1.385 1.665 1.385 1.665 0.605 1.275 0.605 1.275 0.545 1.665 0.545 1.665 0.42 1.545 0.42 1.545 0.36 1.725 0.36 ;
      POLYGON 1.015 0.59 0.335 0.59 0.335 1.09 0.275 1.09 0.275 0.305 0.335 0.305 0.335 0.53 1.015 0.53 ;
  END
END NAND4BBXL

MACRO NAND4BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.623 LAYER Metal1 ;
    ANTENNADIFFAREA 0.8767 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 21.29914525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 161.4358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.84 1.48 0.78 1.48 0.78 1.26 0.42 1.26 0.42 1.48 0.36 1.48 0.36 1.26 0.06 1.26 0.06 0.98 0.08 0.98 0.08 0.44 0.205 0.44 0.205 0.38 0.265 0.38 0.265 0.5 0.14 0.5 0.14 1.2 0.84 1.2 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.76 1.14 1.26 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 0.92 0.65 0.92 0.65 0.43 0.73 0.43 0.73 0.79 0.74 0.79 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.55 1.1 0.47 1.1 0.47 0.92 0.46 0.92 0.46 0.61 0.54 0.61 0.54 0.8 0.55 0.8 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 1.1 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.155 1.65 0.155 1.36 0.215 1.36 0.215 1.65 0.565 1.65 0.565 1.36 0.625 1.36 0.625 1.65 0.985 1.65 0.985 1.36 1.045 1.36 1.045 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 0.97 0.06 0.97 0.5 0.91 0.5 0.91 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.3 1.21 1.24 1.21 1.24 0.66 0.96 0.66 0.96 0.805 0.84 0.805 0.84 0.745 0.9 0.745 0.9 0.6 1.145 0.6 1.145 0.52 1.205 0.52 1.205 0.6 1.3 0.6 ;
  END
END NAND4BX1

MACRO NAND4BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX2 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.337775 LAYER Metal1 ;
    ANTENNADIFFAREA 1.7184 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 22.86794875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 173.69230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.355 0.515 2.28 0.515 2.28 0.715 1.24 0.715 1.24 1.115 2.205 1.115 2.205 1.395 2.115 1.395 2.115 1.175 1.765 1.175 1.765 1.395 1.705 1.395 1.705 1.175 1.355 1.175 1.355 1.395 1.295 1.395 1.295 1.3 1.26 1.3 1.26 1.175 0.945 1.175 0.945 1.395 0.885 1.395 0.885 1.115 1.18 1.115 1.18 0.655 2.22 0.655 2.22 0.455 2.355 0.455 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.42 0.895 0.18 0.895 0.18 0.79 0.03 0.79 0.03 0.705 0.26 0.705 0.26 0.815 0.42 0.815 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.17948725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.34 0.815 1.565 1.015 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.045 1.015 1.665 1.015 1.665 0.815 1.965 0.815 1.965 0.85 2.045 0.85 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.57 0.97 2.145 0.97 2.145 0.89 2.16 0.89 2.16 0.815 2.57 0.815 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 1.77 0 1.77 0 1.65 0.105 1.65 0.105 0.995 0.165 0.995 0.165 1.65 0.68 1.65 0.68 1.275 0.74 1.275 0.74 1.65 1.09 1.65 1.09 1.275 1.15 1.275 1.15 1.65 1.5 1.65 1.5 1.275 1.56 1.275 1.56 1.65 1.91 1.65 1.91 1.275 1.97 1.275 1.97 1.65 2.32 1.65 2.32 1.07 2.38 1.07 2.38 1.65 2.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 0.06 0.845 0.06 0.845 0.375 0.785 0.375 0.785 0.06 0.205 0.06 0.205 0.2 0.145 0.2 0.145 0.06 0 0.06 0 -0.06 2.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.53 0.415 2.47 0.415 2.47 0.355 2.12 0.355 2.12 0.415 2.06 0.415 2.06 0.355 1.725 0.355 1.725 0.375 1.605 0.375 1.605 0.315 1.675 0.315 1.675 0.295 2.53 0.295 ;
      POLYGON 1.945 0.535 1.885 0.535 1.885 0.555 1.195 0.555 1.195 0.505 1.165 0.505 1.165 0.425 1.285 0.425 1.285 0.475 1.825 0.475 1.825 0.455 1.945 0.455 ;
      POLYGON 1.505 0.345 1.385 0.345 1.385 0.325 1.05 0.325 1.05 0.535 0.58 0.535 0.58 0.395 0.64 0.395 0.64 0.475 0.99 0.475 0.99 0.265 1.435 0.265 1.435 0.285 1.505 0.285 ;
      POLYGON 0.8 0.9 0.6 0.9 0.6 1.02 0.52 1.02 0.52 0.715 0.36 0.715 0.36 0.54 0.44 0.54 0.44 0.635 0.6 0.635 0.6 0.82 0.8 0.82 ;
  END
END NAND4BX2

MACRO NAND4BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BX4 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4556 LAYER Metal1 ;
    ANTENNADIFFAREA 3.1243 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 20.98803425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 166.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.03 0.565 3.16 0.565 3.16 0.715 1.54 0.715 1.54 0.995 3.775 0.995 3.775 1.355 3.715 1.355 3.715 1.055 3.365 1.055 3.365 1.355 3.305 1.355 3.305 1.055 2.81 1.055 2.81 1.355 2.75 1.355 2.75 1.055 2.4 1.055 2.4 1.355 2.34 1.355 2.34 1.055 1.99 1.055 1.99 1.355 1.93 1.355 1.93 1.055 1.58 1.055 1.58 1.355 1.52 1.355 1.52 1.11 1.46 1.11 1.46 1.025 1.155 1.025 1.155 1.355 1.095 1.355 1.095 1.025 0.745 1.025 0.745 1.355 0.685 1.355 0.685 0.965 1.48 0.965 1.48 0.655 3.1 0.655 3.1 0.505 3.535 0.505 3.535 0.425 3.595 0.425 3.595 0.505 3.97 0.505 3.97 0.425 4.03 0.425 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.18 1.06 0.1 1.06 0.1 0.73 0.06 0.73 0.06 0.6 0.14 0.6 0.14 0.65 0.18 0.65 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.64 0.815 2.14 0.895 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.38 0.725 3.32 0.725 3.32 0.895 2.45 0.895 2.45 0.835 3.035 0.835 3.035 0.815 3.26 0.815 3.26 0.665 3.38 0.665 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.82051275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.92 0.745 3.765 0.745 3.765 0.895 3.44 0.895 3.44 0.815 3.62 0.815 3.62 0.665 3.92 0.665 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.075 1.65 0.075 1.16 0.135 1.16 0.135 1.65 0.48 1.65 0.48 0.965 0.54 0.965 0.54 1.65 0.89 1.65 0.89 1.235 0.95 1.235 0.95 1.65 1.3 1.65 1.3 1.235 1.36 1.235 1.36 1.65 1.725 1.65 1.725 1.235 1.785 1.235 1.785 1.65 2.135 1.65 2.135 1.235 2.195 1.235 2.195 1.65 2.545 1.65 2.545 1.235 2.605 1.235 2.605 1.65 2.955 1.65 2.955 1.235 3.015 1.235 3.015 1.65 3.51 1.65 3.51 1.235 3.57 1.235 3.57 1.65 3.92 1.65 3.92 0.965 3.98 0.965 3.98 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 1.155 0.06 1.155 0.425 1.095 0.425 1.095 0.06 0.745 0.06 0.745 0.425 0.685 0.425 0.685 0.06 0.135 0.06 0.135 0.5 0.075 0.5 0.075 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.235 0.405 4.175 0.405 4.175 0.245 3.8 0.245 3.8 0.405 3.74 0.405 3.74 0.245 3.39 0.245 3.39 0.405 3.33 0.405 3.33 0.245 2.84 0.245 2.84 0.375 2.72 0.375 2.72 0.245 2.445 0.245 2.445 0.375 2.31 0.375 2.31 0.315 2.385 0.315 2.385 0.185 4.235 0.185 ;
      POLYGON 3.215 0.405 3 0.405 3 0.555 1.56 0.555 1.56 0.535 1.475 0.535 1.475 0.475 1.61 0.475 1.61 0.495 1.915 0.495 1.915 0.435 1.975 0.435 1.975 0.495 2.545 0.495 2.545 0.425 2.605 0.425 2.605 0.495 2.94 0.495 2.94 0.345 3.215 0.345 ;
      POLYGON 2.21 0.395 2.075 0.395 2.075 0.335 1.8 0.335 1.8 0.395 1.68 0.395 1.68 0.335 1.36 0.335 1.36 0.585 0.48 0.585 0.48 0.445 0.54 0.445 0.54 0.525 0.89 0.525 0.89 0.445 0.95 0.445 0.95 0.525 1.3 0.525 1.3 0.275 2.135 0.275 2.135 0.335 2.21 0.335 ;
      POLYGON 1.055 0.745 0.34 0.745 0.34 1.29 0.28 1.29 0.28 0.52 0.34 0.52 0.34 0.685 1.055 0.685 ;
  END
END NAND4BX4

MACRO NAND4BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4BXL 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.612 LAYER Metal1 ;
    ANTENNADIFFAREA 0.73495 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 37.77777775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 281.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.86 1.215 0.56 1.215 0.56 1.12 0.46 1.12 0.46 1.215 0.34 1.215 0.34 1.12 0.08 1.12 0.08 0.54 0.06 0.54 0.06 0.3 0.215 0.3 0.215 0.24 0.275 0.24 0.275 0.36 0.14 0.36 0.14 1.06 0.62 1.06 0.62 1.155 0.86 1.155 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.165 0.895 1.115 0.895 1.115 1.225 1.035 1.225 1.035 0.775 1.165 0.775 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.23 0.74 0.73 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 0.73 0.46 0.73 0.46 0.25 0.54 0.25 0.54 0.6 0.56 0.6 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.46 0.34 0.96 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.165 1.65 0.165 1.22 0.225 1.22 0.225 1.65 0.535 1.65 0.535 1.51 0.595 1.51 0.595 1.65 1.005 1.65 1.005 1.51 1.065 1.51 1.065 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 1.02 0.06 1.02 0.36 0.96 0.36 0.96 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.325 1.245 1.265 1.245 1.265 0.55 0.855 0.55 0.855 0.49 1.265 0.49 1.265 0.385 1.165 0.385 1.165 0.265 1.225 0.265 1.225 0.325 1.325 0.325 ;
  END
END NAND4BXL

MACRO NAND4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4098 LAYER Metal1 ;
    ANTENNADIFFAREA 0.77615 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.08 0.85 1.08 0.85 1.3 0.79 1.3 0.79 1.08 0.43 1.08 0.43 1.3 0.37 1.3 0.37 1.02 1.04 1.02 1.04 0.54 1.1 0.54 1.1 0.79 1.14 0.79 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.34 0.92 0.03 0.92 0.03 0.84 0.23 0.84 0.23 0.65 0.34 0.65 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 0.89 0.48 0.89 0.48 0.54 0.46 0.54 0.46 0.41 0.54 0.41 0.54 0.46 0.56 0.46 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.076923 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.22 0.74 0.83 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.41 0.94 0.91 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.165 1.65 0.165 1.02 0.225 1.02 0.225 1.65 0.575 1.65 0.575 1.18 0.635 1.18 0.635 1.65 1 1.65 1 1.18 1.06 1.18 1.06 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.325 0.06 0.325 0.52 0.265 0.52 0.265 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NAND4X1

MACRO NAND4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X2 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6609 LAYER Metal1 ;
    ANTENNADIFFAREA 1.6934 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.14 1.345 1.79 1.345 1.79 1.405 1.73 1.405 1.73 1.345 1.32 1.345 1.32 1.405 1.26 1.405 1.26 1.345 0.85 1.345 0.85 1.405 0.79 1.405 0.79 1.345 0.38 1.345 0.38 1.405 0.32 1.405 0.32 1.285 2.06 1.285 2.06 0.525 1.185 0.525 1.185 0.505 1.07 0.505 1.07 0.445 1.235 0.445 1.235 0.465 2.12 0.465 2.12 1.17 2.14 1.17 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 12.051282 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 1.185 0.26 1.185 0.26 0.82 0.32 0.82 0.32 1.125 1.86 1.125 1.86 0.82 1.94 0.82 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.17948725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.66 1.025 0.48 1.025 0.48 0.92 0.46 0.92 0.46 0.895 0.42 0.895 0.42 0.835 0.46 0.835 0.46 0.79 0.54 0.79 0.54 0.965 1.6 0.965 1.6 0.845 1.66 0.845 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.3846155 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.395 0.865 0.685 0.865 0.685 0.805 1.335 0.805 1.335 0.705 1.235 0.705 1.235 0.625 1.395 0.625 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.135 0.705 0.86 0.705 0.86 0.4 0.94 0.4 0.94 0.625 1.135 0.625 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.1 1.65 0.1 1.015 0.16 1.015 0.16 1.65 0.525 1.65 0.525 1.49 0.645 1.49 0.645 1.55 0.585 1.55 0.585 1.65 0.995 1.65 0.995 1.49 1.115 1.49 1.115 1.55 1.055 1.55 1.055 1.65 1.465 1.65 1.465 1.49 1.585 1.49 1.585 1.55 1.525 1.55 1.525 1.65 1.99 1.65 1.99 1.49 2.11 1.49 2.11 1.55 2.05 1.55 2.05 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 1.965 0.06 1.965 0.305 2.025 0.305 2.025 0.365 1.905 0.365 1.905 0.06 0.245 0.06 0.245 0.395 0.185 0.395 0.185 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NAND4X2

MACRO NAND4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X4 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.22005 LAYER Metal1 ;
    ANTENNADIFFAREA 2.90415 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.695 0.585 2.805 0.585 2.805 0.715 1.14 0.715 1.14 0.995 3.44 0.995 3.44 1.365 3.38 1.365 3.38 1.055 3.03 1.055 3.03 1.365 2.97 1.365 2.97 1.055 2.455 1.055 2.455 1.365 2.395 1.365 2.395 1.055 2.045 1.055 2.045 1.365 1.985 1.365 1.985 1.055 1.6 1.055 1.6 1.365 1.54 1.365 1.54 1.055 1.19 1.055 1.19 1.365 1.13 1.365 1.13 1.11 1.06 1.11 1.06 1.035 0.755 1.035 0.755 1.365 0.695 1.365 0.695 1.035 0.335 1.035 0.335 1.365 0.275 1.365 0.275 0.975 1.08 0.975 1.08 0.655 2.745 0.655 2.745 0.525 3.205 0.525 3.205 0.445 3.265 0.445 3.265 0.525 3.635 0.525 3.635 0.445 3.695 0.445 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.23 0.625 0.73 0.705 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.24 0.815 1.74 0.895 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.923077 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.025 0.745 2.965 0.745 2.965 0.895 2.095 0.895 2.095 0.835 2.835 0.835 2.835 0.815 2.905 0.815 2.905 0.685 3.025 0.685 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.76923075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.585 0.765 3.545 0.765 3.545 0.895 3.105 0.895 3.105 0.815 3.465 0.815 3.465 0.685 3.585 0.685 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.975 0.13 0.975 0.13 1.65 0.48 1.65 0.48 1.245 0.54 1.245 0.54 1.65 0.9 1.65 0.9 1.245 0.96 1.245 0.96 1.65 1.335 1.65 1.335 1.245 1.395 1.245 1.395 1.65 1.745 1.65 1.745 1.245 1.805 1.245 1.805 1.65 2.19 1.65 2.19 1.245 2.25 1.245 2.25 1.65 2.6 1.65 2.6 1.245 2.66 1.245 2.66 1.65 3.175 1.65 3.175 1.245 3.235 1.245 3.235 1.65 3.645 1.65 3.645 0.975 3.705 0.975 3.705 1.65 4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 0.775 0.06 0.775 0.365 0.715 0.365 0.715 0.06 0.365 0.06 0.365 0.365 0.305 0.365 0.305 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.9 0.425 3.84 0.425 3.84 0.265 3.47 0.265 3.47 0.425 3.41 0.425 3.41 0.265 3.06 0.265 3.06 0.425 3 0.425 3 0.265 2.485 0.265 2.485 0.395 2.365 0.395 2.365 0.265 2.09 0.265 2.09 0.395 1.955 0.395 1.955 0.335 2.03 0.335 2.03 0.205 3.9 0.205 ;
      POLYGON 2.885 0.425 2.645 0.425 2.645 0.555 1.17 0.555 1.17 0.475 1.095 0.475 1.095 0.415 1.23 0.415 1.23 0.495 1.535 0.495 1.535 0.385 1.595 0.385 1.595 0.495 2.19 0.495 2.19 0.435 2.25 0.435 2.25 0.495 2.585 0.495 2.585 0.365 2.885 0.365 ;
      POLYGON 1.83 0.335 1.695 0.335 1.695 0.285 1.42 0.285 1.42 0.335 1.3 0.335 1.3 0.285 0.98 0.285 0.98 0.525 0.1 0.525 0.1 0.385 0.16 0.385 0.16 0.465 0.51 0.465 0.51 0.385 0.57 0.385 0.57 0.465 0.92 0.465 0.92 0.225 1.755 0.225 1.755 0.275 1.83 0.275 ;
  END
END NAND4X4

MACRO NAND4X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X6 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6051 LAYER Metal1 ;
    ANTENNADIFFAREA 4.0665 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.74 0.66 4.32 0.66 4.32 0.79 4.34 0.79 4.34 0.92 4.32 0.92 4.32 1.02 4.475 1.02 4.475 0.9 4.535 0.9 4.535 1.37 4.475 1.37 4.475 1.08 4.125 1.08 4.125 1.37 4.065 1.37 4.065 1.15 3.635 1.15 3.635 1.37 3.575 1.37 3.575 1.01 3.225 1.01 3.225 1.37 3.165 1.37 3.165 1.08 2.755 1.08 2.755 1.37 2.695 1.37 2.695 1.08 2.345 1.08 2.345 1.37 2.285 1.37 2.285 1.08 1.86 1.08 1.86 1.37 1.8 1.37 1.8 1.08 1.31 1.08 1.31 1.37 1.25 1.37 1.25 1.15 0.9 1.15 0.9 1.37 0.84 1.37 0.84 1.15 0.49 1.15 0.49 1.37 0.43 1.37 0.43 0.92 0.49 0.92 0.49 1.09 0.84 1.09 0.84 0.9 0.9 0.9 0.9 1.09 1.25 1.09 1.25 0.9 1.31 0.9 1.31 1.02 2.285 1.02 2.285 0.9 2.345 0.9 2.345 1.02 2.695 1.02 2.695 0.92 2.755 0.92 2.755 1.02 3.165 1.02 3.165 0.95 3.575 0.95 3.575 0.9 3.635 0.9 3.635 1.09 4.065 1.09 4.065 0.92 4.125 0.92 4.125 1.02 4.26 1.02 4.26 0.64 3.825 0.64 3.825 0.52 3.885 0.52 3.885 0.58 4.26 0.58 4.26 0.52 4.32 0.52 4.32 0.6 4.68 0.6 4.68 0.35 4.74 0.35 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 0.991453 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 0.965 0.66 0.965 0.66 0.82 0.385 0.82 0.385 0.74 0.74 0.74 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 0.991453 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.06 0.85 1.74 0.85 1.74 0.92 1.66 0.92 1.66 0.74 1.74 0.74 1.74 0.77 2.06 0.77 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 0.991453 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.095 0.85 2.94 0.85 2.94 0.92 2.86 0.92 2.86 0.85 2.835 0.85 2.835 0.82 2.735 0.82 2.735 0.74 2.915 0.74 2.915 0.77 3.015 0.77 3.015 0.73 3.095 0.73 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 0.991453 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.16 0.82 3.965 0.82 3.965 0.895 3.735 0.895 3.735 0.815 3.86 0.815 3.86 0.74 4.16 0.74 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 1.77 0 1.77 0 1.65 0.225 1.65 0.225 0.9 0.285 0.9 0.285 1.65 0.635 1.65 0.635 1.25 0.695 1.25 0.695 1.65 1.045 1.65 1.045 1.25 1.105 1.25 1.105 1.65 1.595 1.65 1.595 1.25 1.655 1.25 1.655 1.65 2.08 1.65 2.08 1.25 2.14 1.25 2.14 1.65 2.49 1.65 2.49 1.25 2.55 1.25 2.55 1.65 2.9 1.65 2.9 1.25 2.96 1.25 2.96 1.65 3.37 1.65 3.37 1.25 3.43 1.25 3.43 1.65 3.825 1.65 3.825 1.25 3.885 1.25 3.885 1.65 4.27 1.65 4.27 1.25 4.33 1.25 4.33 1.65 4.68 1.65 4.68 0.9 4.74 0.9 4.74 1.65 5 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 0.06 1.105 0.06 1.105 0.47 1.045 0.47 1.045 0.06 0.695 0.06 0.695 0.47 0.635 0.47 0.635 0.06 0.285 0.06 0.285 0.66 0.225 0.66 0.225 0.06 0 0.06 0 -0.06 5 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.535 0.47 4.475 0.47 4.475 0.41 4.09 0.41 4.09 0.47 4.03 0.47 4.03 0.41 3.635 0.41 3.635 0.66 3.575 0.66 3.575 0.41 3.17 0.41 3.17 0.47 3.11 0.47 3.11 0.41 2.76 0.41 2.76 0.47 2.7 0.47 2.7 0.35 4.535 0.35 ;
      POLYGON 3.375 0.63 2.415 0.63 2.415 0.41 2.065 0.41 2.065 0.47 2.005 0.47 2.005 0.41 1.655 0.41 1.655 0.47 1.595 0.47 1.595 0.35 2.475 0.35 2.475 0.57 2.905 0.57 2.905 0.51 2.965 0.51 2.965 0.57 3.315 0.57 3.315 0.51 3.375 0.51 ;
      POLYGON 2.27 0.64 0.43 0.64 0.43 0.35 0.49 0.35 0.49 0.58 0.84 0.58 0.84 0.35 0.9 0.35 0.9 0.58 1.25 0.58 1.25 0.35 1.31 0.35 1.31 0.58 1.8 0.58 1.8 0.52 1.86 0.52 1.86 0.58 2.21 0.58 2.21 0.52 2.27 0.52 ;
  END
END NAND4X6

MACRO NAND4X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4X8 0 0 ;
  SIZE 6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.13415 LAYER Metal1 ;
    ANTENNADIFFAREA 4.844 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.915 0.63 5.54 0.63 5.54 0.73 5.52 0.73 5.52 0.995 5.62 0.995 5.62 0.945 5.68 0.945 5.68 1.39 5.62 1.39 5.62 1.055 5.27 1.055 5.27 1.39 5.21 1.39 5.21 1.08 4.86 1.08 4.86 1.39 4.8 1.39 4.8 1.08 4.45 1.08 4.45 1.39 4.39 1.39 4.39 1.08 4.04 1.08 4.04 1.39 3.98 1.39 3.98 1.08 3.63 1.08 3.63 1.39 3.57 1.39 3.57 1.08 3.22 1.08 3.22 1.39 3.16 1.39 3.16 1.03 2.81 1.03 2.81 1.39 2.75 1.39 2.75 1.03 2.4 1.03 2.4 1.39 2.34 1.39 2.34 1.08 1.99 1.08 1.99 1.39 1.93 1.39 1.93 1.08 1.58 1.08 1.58 1.39 1.52 1.39 1.52 1.08 1.17 1.08 1.17 1.39 1.11 1.39 1.11 1.08 0.76 1.08 0.76 1.39 0.7 1.39 0.7 1.17 0.35 1.17 0.35 1.39 0.29 1.39 0.29 0.97 0.35 0.97 0.35 1.11 0.7 1.11 0.7 0.97 0.76 0.97 0.76 1.02 1.52 1.02 1.52 0.945 1.58 0.945 1.58 1.02 2.34 1.02 2.34 0.97 2.75 0.97 2.75 0.945 2.81 0.945 2.81 0.97 3.16 0.97 3.16 0.945 3.22 0.945 3.22 1.02 3.57 1.02 3.57 0.945 3.63 0.945 3.63 1.02 4.39 1.02 4.39 0.945 4.45 0.945 4.45 1.02 4.8 1.02 4.8 0.995 4.86 0.995 4.86 1.02 5.21 1.02 5.21 0.995 5.46 0.995 5.46 0.63 4.565 0.63 4.565 0.57 5.915 0.57 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 0.984556 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.03 0.905 0.94 0.905 0.94 0.92 0.86 0.92 0.86 0.87 0.4 0.87 0.4 0.79 0.95 0.79 0.95 0.785 1.03 0.785 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 0.984556 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.495 0.87 2.14 0.87 2.14 0.92 2.06 0.92 2.06 0.905 1.865 0.905 1.865 0.785 1.945 0.785 1.945 0.79 2.495 0.79 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.113256 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.94 0.92 3.86 0.92 3.86 0.845 3.27 0.845 3.27 0.785 3.84 0.785 3.84 0.725 3.92 0.725 3.92 0.79 3.94 0.79 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 0.945946 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.705 0.815 5.36 0.895 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 1.77 0 1.77 0 1.65 0.085 1.65 0.085 0.945 0.145 0.945 0.145 1.65 0.495 1.65 0.495 1.27 0.555 1.27 0.555 1.65 0.905 1.65 0.905 1.27 0.965 1.27 0.965 1.65 1.315 1.65 1.315 1.27 1.375 1.27 1.375 1.65 1.725 1.65 1.725 1.27 1.785 1.27 1.785 1.65 2.135 1.65 2.135 1.27 2.195 1.27 2.195 1.65 2.545 1.65 2.545 1.27 2.605 1.27 2.605 1.65 2.955 1.65 2.955 1.27 3.015 1.27 3.015 1.65 3.365 1.65 3.365 1.27 3.425 1.27 3.425 1.65 3.775 1.65 3.775 1.27 3.835 1.27 3.835 1.65 4.185 1.65 4.185 1.27 4.245 1.27 4.245 1.65 4.595 1.65 4.595 1.27 4.655 1.27 4.655 1.65 5.005 1.65 5.005 1.27 5.065 1.27 5.065 1.65 5.415 1.65 5.415 1.27 5.475 1.27 5.475 1.65 5.825 1.65 5.825 0.945 5.885 0.945 5.885 1.65 6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 0.06 1.375 0.06 1.375 0.485 1.315 0.485 1.315 0.06 0.965 0.06 0.965 0.485 0.905 0.485 0.905 0.06 0.555 0.06 0.555 0.485 0.495 0.485 0.495 0.06 0.145 0.06 0.145 0.485 0.085 0.485 0.085 0.06 0 0.06 0 -0.06 6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 3.13 0.395 5.71 0.455 ;
      POLYGON 4.275 0.615 2.955 0.615 2.955 0.47 1.695 0.47 1.695 0.41 3.015 0.41 3.015 0.555 4.275 0.555 ;
      POLYGON 2.84 0.63 2.575 0.63 2.575 0.645 0.35 0.645 0.35 0.63 0.26 0.63 0.26 0.57 0.395 0.57 0.395 0.585 0.67 0.585 0.67 0.57 0.79 0.57 0.79 0.585 1.08 0.585 1.08 0.57 1.2 0.57 1.2 0.585 1.49 0.585 1.49 0.57 1.61 0.57 1.61 0.585 1.9 0.585 1.9 0.57 2.02 0.57 2.02 0.585 2.31 0.585 2.31 0.57 2.43 0.57 2.43 0.585 2.53 0.585 2.53 0.57 2.84 0.57 ;
  END
END NAND4X8

MACRO NAND4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4XL 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3141 LAYER Metal1 ;
    ANTENNADIFFAREA 0.5868 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 1.07 0.86 1.07 0.86 1.05 0.205 1.05 0.205 0.99 0.86 0.99 0.86 0.635 0.845 0.635 0.845 0.515 0.94 0.515 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.1 0.355 0.18 0.855 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.425926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 0.48 0.38 0.855 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.5 0.64 0.58 0.915 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.7 0.64 0.78 0.915 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.285 0.13 1.285 0.13 1.65 0.4 1.65 0.4 1.285 0.46 1.285 0.46 1.65 0.8 1.65 0.8 1.285 0.86 1.285 0.86 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.145 0.06 0.145 0.2 0.085 0.2 0.085 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NAND4XL

MACRO NOR2BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX1 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4236 LAYER Metal1 ;
    ANTENNADIFFAREA 0.51295 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.48205125 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 117.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.32 0.525 0.105 0.525 0.105 0.98 0.185 0.98 0.185 1.455 0.125 1.455 0.125 1.115 0.045 1.115 0.045 0.465 0.26 0.465 0.26 0.355 0.32 0.355 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.575 0.785 0.74 0.945 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.025641 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.365 0.735 0.28 0.735 0.28 0.89 0.165 0.89 0.165 0.6 0.365 0.6 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.77 0 1.77 0 1.65 0.435 1.65 0.435 1.205 0.495 1.205 0.495 1.65 0.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 0.06 0.525 0.06 0.525 0.59 0.465 0.59 0.465 0.06 0.155 0.06 0.155 0.205 0.095 0.205 0.095 0.06 0 0.06 0 -0.06 0.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.73 0.71 0.515 0.71 0.515 1.005 0.73 1.005 0.73 1.185 0.67 1.185 0.67 1.065 0.455 1.065 0.455 0.985 0.33 0.985 0.33 0.925 0.455 0.925 0.455 0.65 0.67 0.65 0.67 0.495 0.73 0.495 ;
  END
END NOR2BX1

MACRO NOR2BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX2 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7686 LAYER Metal1 ;
    ANTENNADIFFAREA 0.926325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.1384615 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 101.84615375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.05 0.52 0.98 0.52 0.98 0.54 0.14 0.54 0.14 0.86 0.76 0.86 0.76 1.36 0.7 1.36 0.7 0.92 0.06 0.92 0.06 0.79 0.08 0.79 0.08 0.48 0.49 0.48 0.49 0.46 0.61 0.46 0.61 0.48 0.93 0.48 0.93 0.46 1.05 0.46 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.3 1.06 1.14 1.06 1.14 1.14 1.06 1.14 1.06 0.98 1.22 0.98 1.22 0.8 1.3 0.8 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.8 0.94 1.3 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.39 1.65 0.39 1.02 0.45 1.02 0.45 1.65 1.11 1.65 1.11 1.24 1.17 1.24 1.17 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.225 0.06 1.225 0.525 1.165 0.525 1.165 0.06 0.77 0.06 0.77 0.32 0.83 0.32 0.83 0.38 0.71 0.38 0.71 0.06 0.33 0.06 0.33 0.32 0.39 0.32 0.39 0.38 0.27 0.38 0.27 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.46 1.09 1.4 1.09 1.4 0.7 0.425 0.7 0.425 0.64 1.4 0.64 1.4 0.43 1.46 0.43 ;
  END
END NOR2BX2

MACRO NOR2BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BX4 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.112 LAYER Metal1 ;
    ANTENNADIFFAREA 1.4257 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.5042735 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 74.17948725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.565 0.55 0.095 0.55 0.095 0.815 0.165 0.815 0.165 0.895 0.095 0.895 0.095 0.995 1.215 0.995 1.215 1.36 1.155 1.36 1.155 1.055 0.595 1.055 0.595 1.36 0.535 1.36 0.535 1.055 0.035 1.055 0.035 0.49 0.275 0.49 0.275 0.43 0.335 0.43 0.335 0.49 0.685 0.49 0.685 0.43 0.745 0.43 0.745 0.49 1.095 0.49 1.095 0.43 1.155 0.43 1.155 0.49 1.505 0.49 1.505 0.43 1.565 0.43 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.923077 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.58 0.815 1.25 0.895 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.29629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.77 1.06 1.54 1.06 1.54 1.11 1.46 1.11 1.46 0.98 1.69 0.98 1.69 0.81 1.77 0.81 ;
    END
  END AN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.17 1.65 0.17 1.24 0.23 1.24 0.23 1.65 0.845 1.65 0.845 1.24 0.905 1.24 0.905 1.65 1.615 1.65 1.615 1.24 1.675 1.24 1.675 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 1.77 0.06 1.77 0.535 1.71 0.535 1.71 0.06 1.33 0.06 1.33 0.33 1.39 0.33 1.39 0.39 1.27 0.39 1.27 0.06 0.92 0.06 0.92 0.33 0.98 0.33 0.98 0.39 0.86 0.39 0.86 0.06 0.51 0.06 0.51 0.33 0.57 0.33 0.57 0.39 0.45 0.39 0.45 0.06 0.1 0.06 0.1 0.33 0.16 0.33 0.16 0.39 0.04 0.39 0.04 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.975 0.56 1.93 0.56 1.93 1.09 1.87 1.09 1.87 0.71 0.905 0.71 0.905 0.715 0.785 0.715 0.785 0.71 0.205 0.71 0.205 0.65 1.87 0.65 1.87 0.5 1.915 0.5 1.915 0.44 1.975 0.44 ;
  END
END NOR2BX4

MACRO NOR2BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2BXL 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4718 LAYER Metal1 ;
    ANTENNADIFFAREA 0.4345 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 29.12345675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 229.62962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.395 0.54 0.14 0.54 0.14 1.24 0.29 1.24 0.29 1.36 0.23 1.36 0.23 1.3 0.06 1.3 0.06 1.17 0.08 1.17 0.08 0.48 0.335 0.48 0.335 0.285 0.395 0.285 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.645 1.06 0.54 1.06 0.54 1.11 0.46 1.11 0.46 0.98 0.565 0.98 0.565 0.715 0.645 0.715 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.64 0.34 1.14 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.54 1.65 0.54 1.24 0.6 1.24 0.6 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.6 0.06 0.6 0.38 0.54 0.38 0.54 0.06 0.19 0.06 0.19 0.38 0.13 0.38 0.13 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.805 1.265 0.745 1.265 0.745 0.6 0.495 0.6 0.495 0.48 0.555 0.48 0.555 0.54 0.745 0.54 0.745 0.285 0.805 0.285 ;
  END
END NOR2BXL

MACRO NOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X1 0 0 ;
  SIZE 0.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2367 LAYER Metal1 ;
    ANTENNADIFFAREA 0.43045 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.515 0.73 0.495 0.73 0.495 1.29 0.435 1.29 0.435 0.65 0.275 0.65 0.275 0.35 0.335 0.35 0.335 0.59 0.515 0.59 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.12820525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.075 0.665 0.195 0.85 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.375 1.085 0.275 1.085 0.275 1.005 0.295 1.005 0.295 0.73 0.375 0.73 ;
    END
  END B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 0.06 0.54 0.06 0.54 0.2 0.42 0.2 0.42 0.06 0.13 0.06 0.13 0.59 0.07 0.59 0.07 0.06 0 0.06 0 -0.06 0.6 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.915 0.13 0.915 0.13 1.65 0.6 1.65 ;
    END
  END VDD
END NOR2X1

MACRO NOR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X2 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3912 LAYER Metal1 ;
    ANTENNADIFFAREA 0.6709 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.955 0.95 0.695 0.95 0.695 1.23 0.54 1.23 0.54 1.41 0.48 1.41 0.48 1.17 0.635 1.17 0.635 0.89 0.895 0.89 0.895 0.73 0.86 0.73 0.86 0.71 0.275 0.71 0.275 0.37 0.335 0.37 0.335 0.65 0.685 0.65 0.685 0.37 0.745 0.37 0.745 0.59 0.955 0.59 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.076923 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.565 1.11 0.38 1.11 0.38 0.89 0.505 0.89 0.505 0.97 0.565 0.97 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.64102575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.815 0.83 0.175 0.83 0.175 0.92 0.06 0.92 0.06 0.77 0.815 0.77 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.94 0.06 0.94 0.2 0.82 0.2 0.82 0.06 0.54 0.06 0.54 0.5 0.48 0.5 0.48 0.06 0.13 0.06 0.13 0.63 0.07 0.63 0.07 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.17 1.65 0.17 1.02 0.23 1.02 0.23 1.65 0.79 1.65 0.79 1.05 0.85 1.05 0.85 1.65 1 1.65 ;
    END
  END VDD
END NOR2X2

MACRO NOR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X4 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6794 LAYER Metal1 ;
    ANTENNADIFFAREA 1.2403 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 0.995 1.44 0.995 1.44 1.125 1.265 1.125 1.265 1.43 1.205 1.43 1.205 1.125 0.6 1.125 0.6 1.43 0.54 1.43 0.54 1.06 1.38 1.06 1.38 0.915 1.675 0.915 1.675 0.73 0.235 0.73 0.235 0.37 0.295 0.37 0.295 0.67 0.645 0.67 0.645 0.37 0.705 0.37 0.705 0.67 1.055 0.67 1.055 0.37 1.115 0.37 1.115 0.67 1.465 0.67 1.465 0.37 1.525 0.37 1.525 0.67 1.74 0.67 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.0897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.285 0.97 1.14 0.97 1.14 0.99 1.06 0.99 1.06 0.97 0.55 0.97 0.55 0.91 1.285 0.91 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.87179475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.595 0.85 0.34 0.85 0.34 0.87 0.26 0.87 0.26 0.85 0.165 0.85 0.165 0.79 1.595 0.79 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.73 0.06 1.73 0.61 1.67 0.61 1.67 0.06 1.32 0.06 1.32 0.61 1.26 0.61 1.26 0.06 0.91 0.06 0.91 0.61 0.85 0.61 0.85 0.06 0.5 0.06 0.5 0.61 0.44 0.61 0.44 0.06 0.17 0.06 0.17 0.2 0.04 0.2 0.04 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.23 1.65 0.23 1.07 0.29 1.07 0.29 1.65 0.85 1.65 0.85 1.19 0.91 1.19 0.91 1.65 1.57 1.65 1.57 1.07 1.63 1.07 1.63 1.65 1.8 1.65 ;
    END
  END VDD
END NOR2X4

MACRO NOR2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X6 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8832 LAYER Metal1 ;
    ANTENNADIFFAREA 1.6883 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.98 0.665 0.125 0.665 0.125 0.905 0.475 0.905 0.475 1.025 1.805 1.025 1.805 1.01 1.885 1.01 1.885 1.395 1.825 1.395 1.825 1.09 1.26 1.09 1.26 1.395 1.2 1.395 1.2 1.09 0.64 1.09 0.64 1.395 0.58 1.395 0.58 1.09 0.415 1.09 0.415 0.965 0.06 0.965 0.06 0.6 0.275 0.6 0.275 0.3 0.335 0.3 0.335 0.6 0.685 0.6 0.685 0.3 0.745 0.3 0.745 0.6 1.095 0.6 1.095 0.3 1.155 0.3 1.155 0.6 1.505 0.6 1.505 0.3 1.565 0.3 1.565 0.6 1.92 0.6 1.92 0.3 1.98 0.3 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.17505 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.46786625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.915 0.905 1.135 0.905 1.135 0.925 1.055 0.925 1.055 0.905 0.555 0.905 0.555 0.845 1.915 0.845 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.17505 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.63324775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.13 0.895 2.07 0.895 2.07 0.785 0.38 0.785 0.38 0.81 0.3 0.81 0.3 0.785 0.205 0.785 0.205 0.725 2.13 0.725 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 0.06 2.185 0.06 2.185 0.54 2.125 0.54 2.125 0.06 1.77 0.06 1.77 0.54 1.71 0.54 1.71 0.06 1.36 0.06 1.36 0.54 1.3 0.54 1.3 0.06 0.95 0.06 0.95 0.54 0.89 0.54 0.89 0.06 0.54 0.06 0.54 0.54 0.48 0.54 0.48 0.06 0.13 0.06 0.13 0.54 0.07 0.54 0.07 0.06 0 0.06 0 -0.06 2.4 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 1.77 0 1.77 0 1.65 0.27 1.65 0.27 1.025 0.33 1.025 0.33 1.65 0.89 1.65 0.89 1.155 0.95 1.155 0.95 1.65 1.515 1.65 1.515 1.155 1.575 1.155 1.575 1.65 2.135 1.65 2.135 1.025 2.195 1.025 2.195 1.65 2.4 1.65 ;
    END
  END VDD
END NOR2X6

MACRO NOR2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X8 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7538 LAYER Metal1 ;
    ANTENNADIFFAREA 2.20955 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.02 1.125 2.955 1.125 2.955 0.665 0.125 0.665 0.125 0.87 0.475 0.87 0.475 1.06 2.77 1.06 2.77 1.045 2.955 1.045 2.955 1.125 2.505 1.125 2.505 1.43 2.445 1.43 2.445 1.125 1.885 1.125 1.885 1.43 1.825 1.43 1.825 1.125 1.26 1.125 1.26 1.43 1.2 1.43 1.2 1.125 0.64 1.125 0.64 1.43 0.58 1.43 0.58 1.125 0.415 1.125 0.415 0.93 0.06 0.93 0.06 0.6 0.275 0.6 0.275 0.3 0.335 0.3 0.335 0.6 0.685 0.6 0.685 0.3 0.745 0.3 0.745 0.6 1.095 0.6 1.095 0.3 1.155 0.3 1.155 0.6 1.505 0.6 1.505 0.3 1.565 0.3 1.565 0.6 1.92 0.6 1.92 0.3 1.98 0.3 1.98 0.6 2.34 0.6 2.34 0.295 2.4 0.295 2.4 0.6 2.75 0.6 2.75 0.3 2.815 0.3 2.815 0.6 3.02 0.6 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.86357775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.7 0.905 1.135 0.905 1.135 0.925 1.055 0.925 1.055 0.905 0.555 0.905 0.555 0.845 2.7 0.845 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.063063 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.5 0.785 0.38 0.785 0.38 0.81 0.3 0.81 0.3 0.785 0.205 0.785 0.205 0.725 2.5 0.725 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 0.06 3.015 0.06 3.015 0.54 2.955 0.54 2.955 0.06 2.605 0.06 2.605 0.54 2.545 0.54 2.545 0.06 2.185 0.06 2.185 0.54 2.125 0.54 2.125 0.06 1.77 0.06 1.77 0.54 1.71 0.54 1.71 0.06 1.36 0.06 1.36 0.54 1.3 0.54 1.3 0.06 0.95 0.06 0.95 0.54 0.89 0.54 0.89 0.06 0.54 0.06 0.54 0.54 0.48 0.54 0.48 0.06 0.13 0.06 0.13 0.54 0.07 0.54 0.07 0.06 0 0.06 0 -0.06 3.2 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 1.77 0 1.77 0 1.65 0.27 1.65 0.27 1.06 0.33 1.06 0.33 1.65 0.89 1.65 0.89 1.19 0.95 1.19 0.95 1.65 1.515 1.65 1.515 1.19 1.575 1.19 1.575 1.65 2.135 1.65 2.135 1.19 2.195 1.19 2.195 1.65 3.2 1.65 ;
    END
  END VDD
END NOR2X8

MACRO NOR2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2XL 0 0 ;
  SIZE 0.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2088 LAYER Metal1 ;
    ANTENNADIFFAREA 0.3523 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.525 1.145 0.435 1.145 0.435 1.005 0.465 1.005 0.465 0.625 0.27 0.625 0.27 0.505 0.33 0.505 0.33 0.565 0.525 0.565 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.17 0.81 0.07 0.81 0.07 0.73 0.08 0.73 0.08 0.545 0.17 0.545 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.4074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.405 0.89 0.35 0.89 0.35 0.97 0.27 0.97 0.27 0.825 0.34 0.825 0.34 0.705 0.405 0.705 ;
    END
  END B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 0.06 0.495 0.06 0.495 0.335 0.435 0.335 0.435 0.06 0.165 0.06 0.165 0.335 0.105 0.335 0.105 0.06 0 0.06 0 -0.06 0.6 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 1.77 0 1.77 0 1.65 0.125 1.65 0.125 1.12 0.185 1.12 0.185 1.65 0.6 1.65 ;
    END
  END VDD
END NOR2XL

MACRO NOR3BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5713 LAYER Metal1 ;
    ANTENNADIFFAREA 0.70025 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.531624 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 145.5384615 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.69 0.49 0.2 0.49 0.2 0.97 0.305 0.97 0.305 1.33 0.245 1.33 0.245 1.03 0.13 1.03 0.13 0.73 0.12 0.73 0.12 0.6 0.13 0.6 0.13 0.24 0.28 0.24 0.28 0.43 0.63 0.43 0.63 0.24 0.69 0.24 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.945 0.895 0.79 0.895 0.79 0.815 0.825 0.815 0.825 0.73 0.945 0.73 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.5641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.55 0.54 1.11 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.051282 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.27 0.575 0.35 0.89 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.715 1.65 0.715 0.97 0.775 0.97 0.775 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.895 0.06 0.895 0.35 0.835 0.35 0.835 0.06 0.485 0.06 0.485 0.35 0.425 0.35 0.425 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.1 1.06 1.04 1.06 1.04 0.67 0.665 0.67 0.665 0.61 1.04 0.61 1.04 0.255 1.1 0.255 ;
  END
END NOR3BX1

MACRO NOR3BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9524 LAYER Metal1 ;
    ANTENNADIFFAREA 1.3306 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.280342 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 125.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.5 0.38 0.14 0.38 0.14 0.86 0.895 0.86 0.895 1.32 0.835 1.32 0.835 0.92 0.06 0.92 0.06 0.79 0.08 0.79 0.08 0.32 1.5 0.32 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.235 1.06 1.235 1.06 0.88 0.995 0.88 0.995 0.8 1.14 0.8 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.3846155 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.92 1.26 0.92 1.26 0.7 0.57 0.7 0.57 0.64 1.34 0.64 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 0.92 1.68 0.92 1.68 1.08 1.6 1.08 1.6 0.64 1.74 0.64 ;
    END
  END AN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.365 1.65 0.365 1.02 0.425 1.02 0.425 1.65 1.515 1.65 1.515 1.18 1.575 1.18 1.575 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.675 0.06 1.675 0.38 1.615 0.38 1.615 0.06 1.205 0.06 1.205 0.16 1.265 0.16 1.265 0.22 1.145 0.22 1.145 0.06 0.735 0.06 0.735 0.16 0.795 0.16 0.795 0.22 0.675 0.22 0.675 0.06 0.265 0.06 0.265 0.16 0.325 0.16 0.325 0.22 0.205 0.22 0.205 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.9 1.08 1.84 1.08 1.84 1.14 1.78 1.14 1.78 1.02 1.84 1.02 1.84 0.54 1.5 0.54 1.5 0.69 1.44 0.69 1.44 0.54 0.47 0.54 0.47 0.68 0.41 0.68 0.41 0.48 1.84 0.48 1.84 0.285 1.9 0.285 ;
  END
END NOR3BX2

MACRO NOR3BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BX4 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.6214 LAYER Metal1 ;
    ANTENNADIFFAREA 2.5687 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.85811975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 104.64102575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.895 0.435 0.315 0.435 0.315 1.125 2.235 1.125 2.235 1.375 2.175 1.375 2.175 1.185 0.985 1.185 0.985 1.375 0.925 1.375 0.925 1.185 0.255 1.185 0.255 0.47 0.14 0.47 0.14 0.54 0.06 0.54 0.06 0.41 0.255 0.41 0.255 0.375 2.895 0.375 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.82051275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.715 0.745 2.65 0.745 2.65 0.865 1.94 0.865 1.94 0.755 1.565 0.755 1.565 0.865 0.66 0.865 0.66 0.6 0.74 0.6 0.74 0.805 1.505 0.805 1.505 0.695 2 0.695 2 0.805 2.59 0.805 2.59 0.685 2.715 0.685 ;
    END
  END B
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.14 0.79 3.02 0.79 3.02 0.705 2.815 0.705 2.815 0.535 3.1 0.535 3.1 0.71 3.14 0.71 ;
    END
  END AN
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.285 0.705 2.165 0.705 2.165 0.595 1.405 0.595 1.405 0.705 1.035 0.705 1.035 0.625 1.165 0.625 1.165 0.645 1.345 0.645 1.345 0.535 2.225 0.535 2.225 0.645 2.285 0.645 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 1.77 0 1.77 0 1.65 0.32 1.65 0.32 1.285 0.44 1.285 0.44 1.345 0.38 1.345 0.38 1.65 1.525 1.65 1.525 1.285 1.645 1.285 1.645 1.345 1.585 1.345 1.585 1.65 2.91 1.65 2.91 1.05 2.97 1.05 2.97 1.65 3.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 0.06 3.07 0.06 3.07 0.435 3.01 0.435 3.01 0.06 2.6 0.06 2.6 0.16 2.66 0.16 2.66 0.22 2.54 0.22 2.54 0.06 2.13 0.06 2.13 0.16 2.19 0.16 2.19 0.22 2.07 0.22 2.07 0.06 1.66 0.06 1.66 0.16 1.72 0.16 1.72 0.22 1.6 0.22 1.6 0.06 1.19 0.06 1.19 0.16 1.25 0.16 1.25 0.22 1.13 0.22 1.13 0.06 0.72 0.06 0.72 0.16 0.78 0.16 0.78 0.22 0.66 0.22 0.66 0.06 0.25 0.06 0.25 0.16 0.31 0.16 0.31 0.22 0.19 0.22 0.19 0.06 0 0.06 0 -0.06 3.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.36 0.545 3.3 0.545 3.3 0.95 3.175 0.95 3.175 1.375 3.115 1.375 3.115 0.95 2.81 0.95 2.81 1.025 0.415 1.025 0.415 0.825 0.475 0.825 0.475 0.965 1.665 0.965 1.665 0.855 1.785 0.855 1.785 0.965 2.75 0.965 2.75 0.89 2.805 0.89 2.805 0.845 2.925 0.845 2.925 0.89 3.24 0.89 3.24 0.485 3.36 0.485 ;
  END
END NOR3BX4

MACRO NOR3BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3BXL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5654 LAYER Metal1 ;
    ANTENNADIFFAREA 0.54225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 34.9012345 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 272.5925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.64 0.365 0.565 0.365 0.565 0.53 0.14 0.53 0.14 1.23 0.275 1.23 0.275 1.35 0.215 1.35 0.215 1.29 0.08 1.29 0.08 0.73 0.06 0.73 0.06 0.6 0.08 0.6 0.08 0.47 0.14 0.47 0.14 0.275 0.2 0.275 0.2 0.47 0.505 0.47 0.505 0.305 0.64 0.305 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.965 0.895 0.845 0.895 0.845 1.13 0.765 1.13 0.765 0.775 0.825 0.775 0.825 0.75 0.905 0.75 0.905 0.775 0.965 0.775 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.63 0.54 1.13 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.63 0.34 1.13 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.74 1.65 0.74 1.23 0.8 1.23 0.8 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.815 0.06 0.815 0.37 0.755 0.37 0.755 0.06 0.405 0.06 0.405 0.37 0.345 0.37 0.345 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.125 1.195 1.005 1.195 1.005 1.255 0.945 1.255 0.945 1.135 1.065 1.135 1.065 0.555 0.725 0.555 0.725 0.615 0.665 0.615 0.665 0.495 1.065 0.495 1.065 0.395 0.96 0.395 0.96 0.275 1.02 0.275 1.02 0.335 1.125 0.335 ;
  END
END NOR3BXL

MACRO NOR3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X1 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3441 LAYER Metal1 ;
    ANTENNADIFFAREA 0.61635 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 0.715 0.885 0.715 0.885 1.335 0.825 1.335 0.825 0.715 0.45 0.715 0.45 0.35 0.51 0.35 0.51 0.655 0.86 0.655 0.86 0.35 0.92 0.35 0.92 0.575 0.94 0.575 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.076923 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 1.005 0.74 1.005 0.74 1.17 0.66 1.17 0.66 0.775 0.76 0.775 ;
    END
  END C
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.897436 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.34 0.91 0.26 0.91 0.26 0.795 0.215 0.795 0.215 0.715 0.26 0.715 0.26 0.655 0.34 0.655 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.775 0.54 1.085 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.245 1.65 0.245 0.975 0.305 0.975 0.305 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.715 0.06 0.715 0.59 0.655 0.59 0.655 0.06 0.305 0.06 0.305 0.59 0.245 0.59 0.245 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NOR3X1

MACRO NOR3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X2 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5148 LAYER Metal1 ;
    ANTENNADIFFAREA 1.12485 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 0.54 1.52 0.54 1.52 1.08 0.91 1.08 0.91 1.14 0.85 1.14 0.85 1.02 1.46 1.02 1.46 0.38 0.245 0.38 0.245 0.32 1.54 0.32 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.92 0.88 0.565 0.88 0.565 0.895 0.435 0.895 0.435 0.815 0.485 0.815 0.485 0.8 0.92 0.8 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.84615375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.145 0.76 1.14 0.76 1.14 0.92 1.06 0.92 1.06 0.7 0.48 0.7 0.48 0.64 1.145 0.64 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.5641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.315 0.705 1.255 0.705 1.255 0.54 0.14 0.54 0.14 0.73 0.06 0.73 0.06 0.48 1.315 0.48 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.275 1.65 0.275 0.93 0.335 0.93 0.335 1.65 1.29 1.65 1.29 1.23 1.41 1.23 1.41 1.29 1.35 1.29 1.35 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.48 0.06 1.48 0.16 1.54 0.16 1.54 0.22 1.42 0.22 1.42 0.06 1.01 0.06 1.01 0.16 1.07 0.16 1.07 0.22 0.95 0.22 0.95 0.06 0.54 0.06 0.54 0.16 0.6 0.16 0.6 0.22 0.48 0.22 0.48 0.06 0.13 0.06 0.13 0.38 0.07 0.38 0.07 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NOR3X2

MACRO NOR3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X4 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9063 LAYER Metal1 ;
    ANTENNADIFFAREA 2.2662 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.94 0.54 2.92 0.54 2.92 1.185 2.225 1.185 2.225 1.375 2.165 1.375 2.165 1.185 0.975 1.185 0.975 1.375 0.915 1.375 0.915 1.125 2.86 1.125 2.86 0.435 0.255 0.435 0.255 0.375 2.92 0.375 2.92 0.41 2.94 0.41 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.0128205 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.7 1.025 0.515 1.025 0.515 1.01 0.08 1.01 0.08 0.92 0.06 0.92 0.06 0.79 0.14 0.79 0.14 0.95 0.575 0.95 0.575 0.965 1.525 0.965 1.525 0.855 1.645 0.855 1.645 0.965 2.64 0.965 2.64 0.825 2.7 0.825 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.4615385 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.54 0.79 2.47 0.79 2.47 0.73 2.37 0.73 2.37 0.82 1.77 0.82 1.77 0.755 1.425 0.755 1.425 0.865 0.675 0.865 0.675 0.85 0.49 0.85 0.49 0.79 0.735 0.79 0.735 0.805 1.365 0.805 1.365 0.695 1.83 0.695 1.83 0.76 2.31 0.76 2.31 0.67 2.46 0.67 2.46 0.6 2.54 0.6 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.8846155 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.115 0.66 1.995 0.66 1.995 0.595 0.985 0.595 0.985 0.705 0.835 0.705 0.835 0.625 0.925 0.625 0.925 0.535 2.055 0.535 2.055 0.6 2.115 0.6 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.77 0 1.77 0 1.65 0.285 1.65 0.285 1.11 0.345 1.11 0.345 1.65 1.46 1.65 1.46 1.285 1.58 1.285 1.58 1.345 1.52 1.345 1.52 1.65 2.675 1.65 2.675 1.285 2.795 1.285 2.795 1.345 2.735 1.345 2.735 1.65 3 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 0.06 2.9 0.06 2.9 0.225 2.96 0.225 2.96 0.285 2.84 0.285 2.84 0.06 2.43 0.06 2.43 0.16 2.49 0.16 2.49 0.22 2.37 0.22 2.37 0.06 1.96 0.06 1.96 0.16 2.02 0.16 2.02 0.22 1.9 0.22 1.9 0.06 1.49 0.06 1.49 0.16 1.55 0.16 1.55 0.22 1.43 0.22 1.43 0.06 1.02 0.06 1.02 0.16 1.08 0.16 1.08 0.22 0.96 0.22 0.96 0.06 0.55 0.06 0.55 0.16 0.61 0.16 0.61 0.22 0.49 0.22 0.49 0.06 0.14 0.06 0.14 0.39 0.08 0.39 0.08 0.06 0 0.06 0 -0.06 3 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NOR3X4

MACRO NOR3X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X6 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2339 LAYER Metal1 ;
    ANTENNADIFFAREA 3.2829 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.14 1.215 3.595 1.215 3.595 1.275 3.535 1.275 3.535 1.215 2.505 1.215 2.505 1.275 2.445 1.275 2.445 1.215 1.095 1.215 1.095 1.275 1.035 1.275 1.035 1.155 4.06 1.155 4.06 0.98 4.08 0.98 4.08 0.605 3.695 0.605 3.695 0.415 2.345 0.415 2.345 0.575 2.285 0.575 2.285 0.415 0.935 0.415 0.935 0.605 0.405 0.605 0.405 0.295 0.465 0.295 0.465 0.545 0.875 0.545 0.875 0.295 0.935 0.295 0.935 0.355 1.345 0.355 1.345 0.295 1.405 0.295 1.405 0.355 1.815 0.355 1.815 0.295 1.875 0.295 1.875 0.355 2.285 0.355 2.285 0.295 2.345 0.295 2.345 0.355 2.755 0.355 2.755 0.295 2.815 0.295 2.815 0.355 3.225 0.355 3.225 0.295 3.285 0.295 3.285 0.355 3.695 0.355 3.695 0.295 3.755 0.295 3.755 0.545 4.14 0.545 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.17505 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5835475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.965 0.88 3.96 0.88 3.96 1.055 0.33 1.055 0.33 0.895 0.235 0.895 0.235 0.815 0.39 0.815 0.39 0.995 1.585 0.995 1.585 0.885 1.705 0.885 1.705 0.995 2.84 0.995 2.84 0.885 2.96 0.885 2.96 0.995 3.9 0.995 3.9 0.845 3.905 0.845 3.905 0.76 3.965 0.76 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.17505 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.7866325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.795 0.895 3.06 0.895 3.06 0.785 2.74 0.785 2.74 0.895 1.805 0.895 1.805 0.785 1.485 0.785 1.485 0.895 0.505 0.895 0.505 0.835 1.425 0.835 1.425 0.725 1.865 0.725 1.865 0.835 1.965 0.835 1.965 0.775 2.025 0.775 2.025 0.835 2.68 0.835 2.68 0.725 3.12 0.725 3.12 0.835 3.635 0.835 3.635 0.815 3.735 0.815 3.735 0.725 3.795 0.725 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.17505 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.227078 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.565 0.735 3.22 0.735 3.22 0.625 2.58 0.625 2.58 0.735 2.125 0.735 2.125 0.625 1.325 0.625 1.325 0.705 1.155 0.705 1.155 0.735 1.035 0.735 1.035 0.625 1.165 0.625 1.165 0.645 1.265 0.645 1.265 0.565 2.185 0.565 2.185 0.675 2.52 0.675 2.52 0.565 3.28 0.565 3.28 0.675 3.565 0.675 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 1.77 0 1.77 0 1.65 0.3 1.65 0.3 1.155 0.36 1.155 0.36 1.65 1.52 1.65 1.52 1.315 1.64 1.315 1.64 1.375 1.58 1.375 1.58 1.65 2.98 1.65 2.98 1.315 3.1 1.315 3.1 1.375 3.04 1.375 3.04 1.65 3.95 1.65 3.95 1.315 4.07 1.315 4.07 1.375 4.01 1.375 4.01 1.65 4.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 0.06 3.49 0.06 3.49 0.16 3.55 0.16 3.55 0.22 3.43 0.22 3.43 0.06 3.02 0.06 3.02 0.16 3.08 0.16 3.08 0.22 2.96 0.22 2.96 0.06 2.55 0.06 2.55 0.16 2.61 0.16 2.61 0.22 2.49 0.22 2.49 0.06 2.08 0.06 2.08 0.16 2.14 0.16 2.14 0.22 2.02 0.22 2.02 0.06 1.61 0.06 1.61 0.16 1.67 0.16 1.67 0.22 1.55 0.22 1.55 0.06 1.14 0.06 1.14 0.16 1.2 0.16 1.2 0.22 1.08 0.22 1.08 0.06 0.67 0.06 0.67 0.16 0.73 0.16 0.73 0.22 0.61 0.22 0.61 0.06 0.26 0.06 0.26 0.605 0.2 0.605 0.2 0.06 0 0.06 0 -0.06 4.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NOR3X6

MACRO NOR3X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3X8 0 0 ;
  SIZE 5.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5195 LAYER Metal1 ;
    ANTENNADIFFAREA 4.3735 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.165 1.085 4.97 1.085 4.97 1.345 4.91 1.345 4.91 1.15 3.825 1.15 3.825 1.21 3.765 1.21 3.765 1.15 2.31 1.15 2.31 1.21 2.25 1.21 2.25 1.15 1.06 1.15 1.06 1.21 1 1.21 1 1.09 4.91 1.09 4.91 0.9 5.025 0.9 5.025 0.335 0.34 0.335 0.34 0.275 5.16 0.275 5.16 0.335 5.085 0.335 5.085 1.005 5.165 1.005 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.35135125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.31 0.83 4.25 0.83 4.25 0.99 0.515 0.99 0.515 0.895 0.235 0.895 0.235 0.815 0.31 0.815 0.31 0.73 0.37 0.73 0.37 0.835 0.575 0.835 0.575 0.93 1.685 0.93 1.685 0.83 1.625 0.83 1.625 0.77 1.745 0.77 1.745 0.93 2.83 0.93 2.83 0.77 2.95 0.77 2.95 0.83 2.89 0.83 2.89 0.93 4.19 0.93 4.19 0.77 4.31 0.77 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.879022 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.765 0.705 4.635 0.705 4.635 0.685 4.41 0.685 4.41 0.67 4.09 0.67 4.09 0.68 3.975 0.68 3.975 0.83 3.535 0.83 3.535 0.68 3.235 0.68 3.235 0.67 2.68 0.67 2.68 0.68 2.62 0.68 2.62 0.83 2.125 0.83 2.125 0.67 1.97 0.67 1.97 0.73 1.91 0.73 1.91 0.67 1.325 0.67 1.325 0.68 1.265 0.68 1.265 0.83 0.675 0.83 0.675 0.735 0.47 0.735 0.47 0.675 0.735 0.675 0.735 0.77 1.205 0.77 1.205 0.62 1.265 0.62 1.265 0.61 2.185 0.61 2.185 0.77 2.56 0.77 2.56 0.62 2.62 0.62 2.62 0.61 3.295 0.61 3.295 0.62 3.595 0.62 3.595 0.77 3.915 0.77 3.915 0.62 4.03 0.62 4.03 0.61 4.47 0.61 4.47 0.625 4.765 0.625 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.4671815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.925 0.725 4.865 0.725 4.865 0.495 3.755 0.495 3.755 0.61 3.815 0.61 3.815 0.67 3.695 0.67 3.695 0.495 2.405 0.495 2.405 0.67 2.285 0.67 2.285 0.61 2.345 0.61 2.345 0.495 1.07 0.495 1.07 0.67 0.835 0.67 0.835 0.435 4.925 0.435 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.2 1.77 0 1.77 0 1.65 0.265 1.65 0.265 0.995 0.325 0.995 0.325 1.65 1.485 1.65 1.485 1.255 1.605 1.255 1.605 1.315 1.545 1.315 1.545 1.65 2.895 1.65 2.895 1.255 3.015 1.255 3.015 1.315 2.955 1.315 2.955 1.65 4.33 1.65 4.33 1.255 4.45 1.255 4.45 1.315 4.39 1.315 4.39 1.65 5.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.2 0.06 4.925 0.06 4.925 0.17 4.805 0.17 4.805 0.06 4.455 0.06 4.455 0.17 4.335 0.17 4.335 0.06 3.985 0.06 3.985 0.17 3.865 0.17 3.865 0.06 3.515 0.06 3.515 0.17 3.395 0.17 3.395 0.06 3.045 0.06 3.045 0.17 2.925 0.17 2.925 0.06 2.575 0.06 2.575 0.17 2.455 0.17 2.455 0.06 2.105 0.06 2.105 0.17 1.985 0.17 1.985 0.06 1.635 0.06 1.635 0.17 1.515 0.17 1.515 0.06 1.165 0.06 1.165 0.17 1.045 0.17 1.045 0.06 0.695 0.06 0.695 0.17 0.575 0.17 0.575 0.06 0.225 0.06 0.225 0.365 0.165 0.365 0.165 0.06 0 0.06 0 -0.06 5.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NOR3X8

MACRO NOR3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3XL 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3072 LAYER Metal1 ;
    ANTENNADIFFAREA 0.485375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 0.73 0.92 0.73 0.92 1.175 0.9 1.175 0.9 1.235 0.84 1.235 0.84 1.115 0.86 1.115 0.86 0.76 0.405 0.76 0.405 0.505 0.465 0.505 0.465 0.7 0.86 0.7 0.86 0.505 0.94 0.505 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.745 1.015 0.74 1.015 0.74 1.355 0.66 1.355 0.66 0.935 0.665 0.935 0.665 0.86 0.745 0.86 ;
    END
  END C
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.36 1.11 0.03 1.11 0.03 0.86 0.11 0.86 0.11 0.955 0.36 0.955 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.945 0.54 1.445 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.235 1.65 0.235 1.21 0.295 1.21 0.295 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.67 0.06 0.67 0.6 0.61 0.6 0.61 0.06 0.3 0.06 0.3 0.2 0.24 0.2 0.24 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NOR3XL

MACRO NOR4BBX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX1 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8257 LAYER Metal1 ;
    ANTENNADIFFAREA 1.0967 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.11453 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 111.74358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.11 1.095 1.11 1.095 1.405 0.5 1.405 0.5 1.465 0.44 1.465 0.44 1.19 0.5 1.19 0.5 1.345 1.035 1.345 1.035 0.565 0.6 0.565 0.6 0.305 0.66 0.305 0.66 0.505 1.035 0.505 1.035 0.305 1.095 0.305 1.095 0.98 1.14 0.98 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.565 0.925 0.54 0.925 0.54 1.13 0.435 1.13 0.435 0.805 0.565 0.805 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.4615385 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.805 0.755 1.145 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 0.97 1.435 0.97 1.435 0.905 1.365 0.905 1.365 0.785 1.54 0.785 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.72222225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.055 0.69 0.14 1.13 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.285 0.13 1.285 0.13 1.65 1.195 1.65 1.195 1.195 1.255 1.195 1.255 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.315 0.06 1.315 0.53 1.255 0.53 1.255 0.06 0.88 0.06 0.88 0.42 0.82 0.42 0.82 0.06 0.425 0.06 0.425 0.295 0.365 0.295 0.365 0.06 0.13 0.06 0.13 0.33 0.07 0.33 0.07 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.52 0.695 1.265 0.695 1.265 1.045 1.52 1.045 1.52 1.29 1.46 1.29 1.46 1.105 1.2 1.105 1.2 0.695 1.16 0.695 1.16 0.635 1.46 0.635 1.46 0.435 1.52 0.435 ;
      POLYGON 0.935 0.745 0.295 0.745 0.295 1.02 0.235 1.02 0.235 0.54 0.295 0.54 0.295 0.685 0.935 0.685 ;
  END
END NOR4BBX1

MACRO NOR4BBX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX2 0 0 ;
  SIZE 3 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5225 LAYER Metal1 ;
    ANTENNADIFFAREA 1.905075 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.0128205 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 102.051282 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.74 0.73 2.72 0.73 2.72 0.865 2.695 0.865 2.695 1.145 2.635 1.145 2.635 0.805 2.66 0.805 2.66 0.51 1.715 0.51 1.715 0.48 1.33 0.48 1.33 0.46 1.26 0.46 1.26 0.4 1.38 0.4 1.38 0.42 1.715 0.42 1.715 0.36 1.775 0.36 1.775 0.45 2.125 0.45 2.125 0.37 2.185 0.37 2.185 0.45 2.535 0.45 2.535 0.37 2.595 0.37 2.595 0.45 2.72 0.45 2.72 0.6 2.74 0.6 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.56 0.73 2.365 0.73 2.365 0.895 2.225 0.895 2.225 0.65 2.56 0.65 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.125 0.925 1.86 0.925 1.86 0.755 2.045 0.755 2.045 0.61 2.125 0.61 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.595 1.085 0.295 1.085 0.295 1.005 0.515 1.005 0.515 0.805 0.595 0.805 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.595 0.705 0.375 0.705 0.375 0.905 0.295 0.905 0.295 0.625 0.595 0.625 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.77 0 1.77 0 1.65 0.4 1.65 0.4 1.185 0.46 1.185 0.46 1.65 1.1 1.65 1.1 1.075 1.16 1.075 1.16 1.65 3 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 0.06 2.8 0.06 2.8 0.35 2.74 0.35 2.74 0.06 2.39 0.06 2.39 0.35 2.33 0.35 2.33 0.06 1.98 0.06 1.98 0.35 1.92 0.35 1.92 0.06 1.54 0.06 1.54 0.26 1.6 0.26 1.6 0.32 1.48 0.32 1.48 0.06 1.145 0.06 1.145 0.35 1.085 0.35 1.085 0.06 0.46 0.06 0.46 0.365 0.4 0.365 0.4 0.06 0 0.06 0 -0.06 3 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.9 1.305 2.02 1.305 2.02 1.185 2.08 1.185 2.08 1.245 2.43 1.245 2.43 0.995 2.49 0.995 2.49 1.245 2.84 1.245 2.84 0.915 2.9 0.915 ;
      POLYGON 2.285 1.145 2.225 1.145 2.225 1.085 1.57 1.085 1.57 1.145 1.51 1.145 1.51 1.025 2.225 1.025 2.225 0.995 2.285 0.995 ;
      POLYGON 1.775 1.305 1.305 1.305 1.305 0.975 0.955 0.975 0.955 1.305 0.895 1.305 0.895 0.915 1.365 0.915 1.365 1.245 1.715 1.245 1.715 1.185 1.775 1.185 ;
      POLYGON 1.675 0.81 1.365 0.81 1.365 0.64 1.1 0.64 1.1 0.51 0.925 0.51 0.925 0.33 0.62 0.33 0.62 0.525 0.195 0.525 0.195 1.095 0.135 1.095 0.135 0.405 0.225 0.405 0.225 0.465 0.56 0.465 0.56 0.27 0.985 0.27 0.985 0.45 1.16 0.45 1.16 0.58 1.425 0.58 1.425 0.75 1.675 0.75 ;
      POLYGON 1.265 0.8 0.78 0.8 0.78 1.095 0.695 1.095 0.695 0.975 0.72 0.975 0.72 0.43 0.78 0.43 0.78 0.74 1.265 0.74 ;
  END
END NOR4BBX2

MACRO NOR4BBX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBX4 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.458875 LAYER Metal1 ;
    ANTENNADIFFAREA 3.236 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.234 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.50801275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 78.923077 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.31 1.3 4.25 1.3 4.25 1.04 3.94 1.04 3.94 1.11 3.9 1.11 3.9 1.3 3.84 1.3 3.84 0.48 1.255 0.48 1.255 0.36 1.315 0.36 1.315 0.42 1.665 0.42 1.665 0.36 1.725 0.36 1.725 0.42 2.075 0.42 2.075 0.36 2.135 0.36 2.135 0.42 2.485 0.42 2.485 0.36 2.545 0.36 2.545 0.42 2.925 0.42 2.925 0.36 2.985 0.36 2.985 0.42 3.335 0.42 3.335 0.36 3.395 0.36 3.395 0.42 3.775 0.42 3.775 0.36 3.835 0.36 3.835 0.42 3.9 0.42 3.9 0.45 4.185 0.45 4.185 0.37 4.245 0.37 4.245 0.51 3.9 0.51 3.9 0.98 4.31 0.98 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.66 0.61 3.74 1.11 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.86 0.58 2.94 1.08 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.76 0.54 1.26 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.76 0.34 1.26 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.77 0 1.77 0 1.65 0.405 1.65 0.405 1.36 0.465 1.36 0.465 1.65 1.18 1.65 1.18 1.34 1.24 1.34 1.24 1.65 1.59 1.65 1.59 1.23 1.65 1.23 1.65 1.65 4.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 0.06 4.45 0.06 4.45 0.35 4.39 0.35 4.39 0.06 4.04 0.06 4.04 0.35 3.98 0.35 3.98 0.06 3.63 0.06 3.63 0.32 3.51 0.32 3.51 0.06 3.22 0.06 3.22 0.32 3.1 0.32 3.1 0.06 2.78 0.06 2.78 0.32 2.66 0.32 2.66 0.06 2.37 0.06 2.37 0.32 2.25 0.32 2.25 0.06 1.96 0.06 1.96 0.32 1.84 0.32 1.84 0.06 1.55 0.06 1.55 0.32 1.43 0.32 1.43 0.06 1.11 0.06 1.11 0.35 1.05 0.35 1.05 0.06 0.39 0.06 0.39 0.5 0.33 0.5 0.33 0.06 0 0.06 0 -0.06 4.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.515 1.46 2.815 1.46 2.815 1.34 2.875 1.34 2.875 1.4 3.225 1.4 3.225 1.34 3.285 1.34 3.285 1.4 3.635 1.4 3.635 1.21 3.695 1.21 3.695 1.4 4.045 1.4 4.045 1.14 4.105 1.14 4.105 1.4 4.455 1.4 4.455 1.07 4.515 1.07 ;
      POLYGON 3.49 1.3 3.43 1.3 3.43 1.24 3.08 1.24 3.08 1.3 3.02 1.3 3.02 1.24 2.47 1.24 2.47 1.3 2.41 1.3 2.41 1.24 2.06 1.24 2.06 1.3 2 1.3 2 1.18 3.43 1.18 3.43 1.07 3.49 1.07 ;
      POLYGON 2.675 1.46 1.795 1.46 1.795 1.13 1.445 1.13 1.445 1.46 1.385 1.46 1.385 1.13 1.035 1.13 1.035 1.46 0.975 1.46 0.975 1.07 1.855 1.07 1.855 1.4 2.205 1.4 2.205 1.34 2.265 1.34 2.265 1.4 2.615 1.4 2.615 1.34 2.675 1.34 ;
      POLYGON 2.025 0.64 0.81 0.64 0.81 0.42 0.55 0.42 0.55 0.66 0.16 0.66 0.16 1.36 0.26 1.36 0.26 1.48 0.2 1.48 0.2 1.42 0.1 1.42 0.1 0.605 0.125 0.605 0.125 0.52 0.185 0.52 0.185 0.6 0.49 0.6 0.49 0.36 0.87 0.36 0.87 0.58 2.025 0.58 ;
      POLYGON 1.215 0.965 0.71 0.965 0.71 1.13 0.7 1.13 0.7 1.48 0.64 1.48 0.64 1.09 0.65 1.09 0.65 0.52 0.71 0.52 0.71 0.905 1.215 0.905 ;
  END
END NOR4BBX4

MACRO NOR4BBXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BBXL 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9257 LAYER Metal1 ;
    ANTENNADIFFAREA 0.933775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 28.57098775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 218.9814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.92 1.32 0.92 1.32 1.41 0.74 1.41 0.74 1.35 1.26 1.35 1.26 0.51 0.83 0.51 0.83 0.255 0.89 0.255 0.89 0.45 1.26 0.45 1.26 0.255 1.32 0.255 1.32 0.79 1.34 0.79 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 1.15 0.74 1.15 0.74 1.25 0.66 1.25 0.66 0.98 0.68 0.98 0.68 0.77 0.76 0.77 ;
    END
  END D
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.085 1.12 0.94 1.12 0.94 1.125 0.86 1.125 0.86 0.98 1.005 0.98 1.005 0.77 1.085 0.77 ;
    END
  END C
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.765 0.895 1.715 0.895 1.715 1.155 1.525 1.155 1.525 1.075 1.635 1.075 1.635 0.815 1.765 0.815 ;
    END
  END AN
  PIN BN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.03 0.685 0.4 0.895 ;
    END
  END BN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.275 1.65 0.275 0.995 0.335 0.995 0.335 1.65 1.49 1.65 1.49 1.32 1.55 1.32 1.55 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.55 0.06 1.55 0.35 1.49 0.35 1.49 0.06 1.095 0.06 1.095 0.35 1.035 0.35 1.035 0.06 0.655 0.06 0.655 0.2 0.595 0.2 0.595 0.06 0.3 0.06 0.3 0.2 0.24 0.2 0.24 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.925 1.315 1.665 1.315 1.665 1.255 1.865 1.255 1.865 0.535 1.42 0.535 1.42 0.475 1.865 0.475 1.865 0.375 1.695 0.375 1.695 0.255 1.755 0.255 1.755 0.315 1.925 0.315 ;
      POLYGON 1.16 0.67 0.56 0.67 0.56 1.055 0.54 1.055 0.54 1.115 0.48 1.115 0.48 0.995 0.5 0.995 0.5 0.585 0.405 0.585 0.405 0.465 0.465 0.465 0.465 0.525 0.56 0.525 0.56 0.61 1.16 0.61 ;
  END
END NOR4BBXL

MACRO NOR4BX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6354 LAYER Metal1 ;
    ANTENNADIFFAREA 0.859125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 21.723077 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 165.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 0.55 0.17 0.55 0.17 1.17 0.295 1.17 0.295 1.425 0.235 1.425 0.235 1.23 0.11 1.23 0.11 0.73 0.06 0.73 0.06 0.6 0.11 0.6 0.11 0.49 0.34 0.49 0.34 0.41 0.4 0.41 0.4 0.49 0.765 0.49 0.765 0.38 0.825 0.38 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.22222225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.045 0.635 1.14 0.93 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.102564 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.64 0.755 0.945 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.102564 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.785 0.54 1.105 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 0.715 0.34 0.94 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.925 1.65 0.925 1.035 0.985 1.035 0.985 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 1.03 0.06 1.03 0.39 0.97 0.39 0.97 0.06 0.605 0.06 0.605 0.39 0.545 0.39 0.545 0.06 0.195 0.06 0.195 0.39 0.135 0.39 0.135 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.265 1.08 1.255 1.08 1.255 1.25 1.195 1.25 1.195 1.01 1.205 1.01 1.205 0.55 0.95 0.55 0.95 0.695 0.83 0.695 0.83 0.635 0.89 0.635 0.89 0.49 1.205 0.49 1.205 0.41 1.265 0.41 ;
  END
END NOR4BX1

MACRO NOR4BX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX2 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.33855 LAYER Metal1 ;
    ANTENNADIFFAREA 1.78865 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 22.8811965 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 173.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.52 1.135 2.46 1.135 2.46 1.055 1.295 1.055 1.295 0.92 1.26 0.92 1.26 0.79 1.295 0.79 1.295 0.545 0.985 0.545 0.985 0.405 1.045 0.405 1.045 0.485 1.395 0.485 1.395 0.405 1.455 0.405 1.455 0.485 1.845 0.485 1.845 0.405 1.905 0.405 1.905 0.485 2.255 0.485 2.255 0.405 2.315 0.405 2.315 0.545 1.355 0.545 1.355 0.995 2.52 0.995 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.455 0.87 0.14 0.87 0.14 0.92 0.06 0.92 0.06 0.79 0.36 0.79 0.36 0.735 0.455 0.735 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.77 0.895 1.455 0.895 1.455 0.645 1.535 0.645 1.535 0.815 1.635 0.815 1.635 0.8 1.77 0.8 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.895 1.87 0.895 1.87 0.645 2.035 0.645 2.035 0.815 2.2 0.815 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.64102575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.3 0.645 2.565 0.895 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 1.77 0 1.77 0 1.65 0.15 1.65 0.15 1.02 0.21 1.02 0.21 1.65 0.9 1.65 0.9 1.315 1.02 1.315 1.02 1.375 0.96 1.375 0.96 1.65 2.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 0.06 2.52 0.06 2.52 0.385 2.46 0.385 2.46 0.06 2.11 0.06 2.11 0.385 2.05 0.385 2.05 0.06 1.66 0.06 1.66 0.385 1.6 0.385 1.6 0.06 1.25 0.06 1.25 0.385 1.19 0.385 1.19 0.06 0.81 0.06 0.81 0.2 0.75 0.2 0.75 0.06 0.355 0.06 0.355 0.635 0.295 0.635 0.295 0.06 0 0.06 0 -0.06 2.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.725 1.295 2.255 1.295 2.255 1.215 1.905 1.215 1.905 1.275 1.845 1.275 1.845 1.155 2.315 1.155 2.315 1.235 2.665 1.235 2.665 1.015 2.725 1.015 ;
      POLYGON 2.14 1.375 2.08 1.375 2.08 1.435 1.37 1.435 1.37 1.375 1.31 1.375 1.31 1.315 1.43 1.315 1.43 1.375 2.02 1.375 2.02 1.315 2.14 1.315 ;
      POLYGON 1.605 1.275 1.545 1.275 1.545 1.215 1.195 1.215 1.195 1.405 1.135 1.405 1.135 1.215 0.785 1.215 0.785 1.275 0.725 1.275 0.725 1.155 1.135 1.155 1.135 1.02 1.195 1.02 1.195 1.155 1.605 1.155 ;
      POLYGON 0.945 0.865 0.645 0.865 0.645 1.045 0.565 1.045 0.565 0.54 0.645 0.54 0.645 0.785 0.945 0.785 ;
  END
END NOR4BX2

MACRO NOR4BX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BX4 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2281 LAYER Metal1 ;
    ANTENNADIFFAREA 3.0517 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.04358975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 147.4358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.015 1.135 3.955 1.135 3.955 1.055 3.605 1.055 3.605 1.135 3.545 1.135 3.545 1.055 1.765 1.055 1.765 1.085 1.635 1.085 1.635 0.615 0.88 0.615 0.88 0.475 0.94 0.475 0.94 0.555 1.29 0.555 1.29 0.475 1.35 0.475 1.35 0.555 1.7 0.555 1.7 0.475 1.76 0.475 1.76 0.555 2.11 0.555 2.11 0.475 2.17 0.475 2.17 0.555 2.52 0.555 2.52 0.475 2.58 0.475 2.58 0.555 2.93 0.555 2.93 0.475 2.99 0.475 2.99 0.555 3.34 0.555 3.34 0.475 3.4 0.475 3.4 0.555 3.75 0.555 3.75 0.475 3.81 0.475 3.81 0.615 1.695 0.615 1.695 0.995 4.015 0.995 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.285 0.955 0.205 0.955 0.205 0.73 0.06 0.73 0.06 0.6 0.14 0.6 0.14 0.65 0.285 0.65 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.795 0.815 2.295 0.895 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.8846155 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.15 0.895 2.595 0.895 2.595 0.715 2.675 0.715 2.675 0.815 3.15 0.815 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.8846155 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.97 0.895 3.415 0.895 3.415 0.715 3.495 0.715 3.495 0.815 3.97 0.815 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.145 1.65 0.145 1.055 0.205 1.055 0.205 1.65 0.83 1.65 0.83 1.345 0.95 1.345 0.95 1.405 0.89 1.405 0.89 1.65 1.24 1.65 1.24 1.345 1.36 1.345 1.36 1.405 1.3 1.405 1.3 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 4.015 0.06 4.015 0.455 3.955 0.455 3.955 0.06 3.605 0.06 3.605 0.455 3.545 0.455 3.545 0.06 3.195 0.06 3.195 0.455 3.135 0.455 3.135 0.06 2.785 0.06 2.785 0.455 2.725 0.455 2.725 0.06 2.375 0.06 2.375 0.455 2.315 0.455 2.315 0.06 1.965 0.06 1.965 0.455 1.905 0.455 1.905 0.06 1.555 0.06 1.555 0.455 1.495 0.455 1.495 0.06 1.145 0.06 1.145 0.455 1.085 0.455 1.085 0.06 0.705 0.06 0.705 0.2 0.645 0.2 0.645 0.06 0.205 0.06 0.205 0.5 0.145 0.5 0.145 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.22 1.295 3.34 1.295 3.34 1.215 2.99 1.215 2.99 1.275 2.93 1.275 2.93 1.215 2.58 1.215 2.58 1.275 2.52 1.275 2.52 1.155 3.4 1.155 3.4 1.235 3.75 1.235 3.75 1.175 3.81 1.175 3.81 1.235 4.16 1.235 4.16 1.015 4.22 1.015 ;
      POLYGON 3.225 1.375 3.165 1.375 3.165 1.435 1.725 1.435 1.725 1.405 1.665 1.405 1.665 1.345 1.785 1.345 1.785 1.375 2.085 1.375 2.085 1.345 2.205 1.345 2.205 1.375 2.695 1.375 2.695 1.315 2.815 1.315 2.815 1.375 3.105 1.375 3.105 1.315 3.225 1.315 ;
      POLYGON 2.38 1.275 2.32 1.275 2.32 1.215 1.96 1.215 1.96 1.275 1.9 1.275 1.9 1.245 1.535 1.245 1.535 1.435 1.475 1.435 1.475 1.245 1.125 1.245 1.125 1.435 1.065 1.435 1.065 1.245 0.715 1.245 0.715 1.305 0.655 1.305 0.655 1.185 1.065 1.185 1.065 1.045 1.125 1.045 1.125 1.185 1.475 1.185 1.475 1.045 1.535 1.045 1.535 1.185 1.9 1.185 1.9 1.155 2.38 1.155 ;
      POLYGON 1.285 0.775 0.445 0.775 0.445 1.02 0.385 1.02 0.385 0.52 0.445 0.52 0.445 0.715 1.285 0.715 ;
  END
END NOR4BX4

MACRO NOR4BXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4BXL 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7679 LAYER Metal1 ;
    ANTENNADIFFAREA 0.754275 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 47.4012345 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 353.14814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.105 0.35 1.045 0.35 1.045 0.515 0.14 0.515 0.14 1.02 0.535 1.02 0.535 1.14 0.475 1.14 0.475 1.08 0.08 1.08 0.08 0.73 0.06 0.73 0.06 0.6 0.08 0.6 0.08 0.455 0.605 0.455 0.605 0.26 0.665 0.26 0.665 0.455 0.985 0.455 0.985 0.29 1.105 0.29 ;
    END
  END Y
  PIN AN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.565 0.895 1.265 0.895 1.265 0.815 1.38 0.815 1.38 0.615 1.46 0.615 1.46 0.815 1.565 0.815 ;
    END
  END AN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 0.98 1.06 0.98 1.06 0.87 0.925 0.87 0.925 0.615 1.005 0.615 1.005 0.79 1.14 0.79 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.825 0.775 0.765 0.775 0.765 1.085 0.635 1.085 0.635 1.005 0.685 1.005 0.685 0.695 0.825 0.695 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.535 0.92 0.26 0.92 0.26 0.73 0.455 0.73 0.455 0.615 0.535 0.615 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 1.24 1.65 1.24 1.02 1.3 1.02 1.3 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.3 0.06 1.3 0.355 1.24 0.355 1.24 0.06 0.87 0.06 0.87 0.355 0.81 0.355 0.81 0.06 0.46 0.06 0.46 0.355 0.4 0.355 0.4 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.725 1.055 1.505 1.055 1.505 1.115 1.445 1.115 1.445 0.995 1.665 0.995 1.665 0.515 1.225 0.515 1.225 0.575 1.165 0.575 1.165 0.455 1.445 0.455 1.445 0.26 1.505 0.26 1.505 0.455 1.725 0.455 ;
  END
END NOR4BXL

MACRO NOR4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X1 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3524 LAYER Metal1 ;
    ANTENNADIFFAREA 0.71775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 1.495 0.86 1.495 0.86 0.9 0.865 0.9 0.865 0.61 0.235 0.61 0.235 0.49 0.295 0.49 0.295 0.55 0.655 0.55 0.655 0.49 0.715 0.49 0.715 0.55 0.925 0.55 0.925 0.9 0.94 0.9 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.897436 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.22 0.79 0.03 0.79 0.03 0.6 0.14 0.6 0.14 0.67 0.22 0.67 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.5897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.425 1.11 0.26 1.11 0.26 0.98 0.345 0.98 0.345 0.73 0.425 0.73 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.12820525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.585 1.3 0.46 1.3 0.46 1.17 0.525 1.17 0.525 0.73 0.585 0.73 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.4358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.805 0.85 0.74 0.85 0.74 0.92 0.66 0.92 0.66 0.73 0.805 0.73 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.13 1.65 0.13 0.9 0.19 0.9 0.19 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.92 0.06 0.92 0.47 0.86 0.47 0.86 0.06 0.5 0.06 0.5 0.47 0.44 0.47 0.44 0.06 0.17 0.06 0.17 0.2 0.04 0.2 0.04 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NOR4X1

MACRO NOR4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6228 LAYER Metal1 ;
    ANTENNADIFFAREA 1.38625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 1.345 1.01 1.345 1.01 1.285 1.86 1.285 1.86 1.17 1.88 1.17 1.88 0.525 0.345 0.525 0.345 0.505 0.275 0.505 0.275 0.445 0.395 0.445 0.395 0.465 0.715 0.465 0.715 0.445 0.835 0.445 0.835 0.465 1.155 0.465 1.155 0.445 1.275 0.445 1.275 0.465 1.595 0.465 1.595 0.445 1.715 0.445 1.715 0.465 1.94 0.465 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.025641 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 1.185 0.26 1.185 0.26 0.82 0.32 0.82 0.32 1.125 1.66 1.125 1.66 0.98 1.68 0.98 1.68 0.82 1.74 0.82 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.495 1.025 0.48 1.025 0.48 0.92 0.46 0.92 0.46 0.895 0.42 0.895 0.42 0.835 0.46 0.835 0.46 0.79 0.54 0.79 0.54 0.965 1.435 0.965 1.435 0.845 1.495 0.845 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.565 0.705 1.335 0.705 1.335 0.865 0.64 0.865 0.64 0.805 1.275 0.805 1.275 0.625 1.565 0.625 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.64 0.625 1.14 0.705 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.215 1.65 0.215 1.285 0.275 1.285 0.275 1.65 1.67 1.65 1.67 1.54 1.79 1.54 1.79 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.875 0.06 1.875 0.305 1.935 0.305 1.935 0.365 1.815 0.365 1.815 0.06 1.435 0.06 1.435 0.305 1.495 0.305 1.495 0.365 1.375 0.365 1.375 0.06 0.995 0.06 0.995 0.305 1.055 0.305 1.055 0.365 0.935 0.365 0.935 0.06 0.555 0.06 0.555 0.305 0.615 0.305 0.615 0.365 0.495 0.365 0.495 0.06 0.16 0.06 0.16 0.395 0.1 0.395 0.1 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NOR4X2

MACRO NOR4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X4 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.988 LAYER Metal1 ;
    ANTENNADIFFAREA 2.70275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.52 0.655 1.14 0.655 1.14 0.995 3.465 0.995 3.465 1.135 3.405 1.135 3.405 1.055 3.055 1.055 3.055 1.135 2.995 1.135 2.995 1.055 1.08 1.055 1.08 0.92 1.06 0.92 1.06 0.79 1.08 0.79 1.08 0.655 0.59 0.655 0.59 0.515 0.65 0.515 0.65 0.595 1 0.595 1 0.515 1.06 0.515 1.06 0.595 1.41 0.595 1.41 0.515 1.47 0.515 1.47 0.595 1.82 0.595 1.82 0.515 1.88 0.515 1.88 0.595 2.23 0.595 2.23 0.515 2.29 0.515 2.29 0.595 2.64 0.595 2.64 0.515 2.7 0.515 2.7 0.595 3.05 0.595 3.05 0.515 3.11 0.515 3.11 0.595 3.46 0.595 3.46 0.515 3.52 0.515 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.0128205 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 0.95 0.35 0.95 0.35 0.87 0.86 0.87 0.86 0.755 0.94 0.755 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.80769225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.805 0.895 1.24 0.895 1.24 0.815 1.725 0.815 1.725 0.755 1.805 0.755 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.57 0.895 2.11 0.895 2.11 0.815 2.435 0.815 2.435 0.775 2.57 0.775 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.80769225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.42 0.895 2.835 0.895 2.835 0.815 3.105 0.815 3.105 0.775 3.185 0.775 3.185 0.815 3.42 0.815 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.355 0.395 1.355 0.395 1.415 0.335 1.415 0.335 1.65 0.685 1.65 0.685 1.355 0.805 1.355 0.805 1.415 0.745 1.415 0.745 1.65 3.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 0.06 3.725 0.06 3.725 0.495 3.665 0.495 3.665 0.06 3.315 0.06 3.315 0.495 3.255 0.495 3.255 0.06 2.905 0.06 2.905 0.495 2.845 0.495 2.845 0.06 2.495 0.06 2.495 0.495 2.435 0.495 2.435 0.06 2.085 0.06 2.085 0.495 2.025 0.495 2.025 0.06 1.675 0.06 1.675 0.495 1.615 0.495 1.615 0.06 1.265 0.06 1.265 0.495 1.205 0.495 1.205 0.06 0.855 0.06 0.855 0.495 0.795 0.495 0.795 0.06 0.445 0.06 0.445 0.495 0.385 0.495 0.385 0.06 0 0.06 0 -0.06 3.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.67 1.295 2.79 1.295 2.79 1.215 2.44 1.215 2.44 1.275 2.38 1.275 2.38 1.215 2.03 1.215 2.03 1.275 1.97 1.275 1.97 1.155 2.85 1.155 2.85 1.235 3.2 1.235 3.2 1.175 3.26 1.175 3.26 1.235 3.61 1.235 3.61 1.015 3.67 1.015 ;
      POLYGON 2.675 1.375 2.615 1.375 2.615 1.435 1.16 1.435 1.16 1.415 1.1 1.415 1.1 1.355 1.22 1.355 1.22 1.375 1.51 1.375 1.51 1.355 1.63 1.355 1.63 1.375 2.145 1.375 2.145 1.315 2.265 1.315 2.265 1.375 2.555 1.375 2.555 1.315 2.675 1.315 ;
      POLYGON 1.805 1.275 1.745 1.275 1.745 1.215 1.395 1.215 1.395 1.275 1.335 1.275 1.335 1.215 0.98 1.215 0.98 1.445 0.92 1.445 0.92 1.215 0.57 1.215 0.57 1.445 0.51 1.445 0.51 1.255 0.16 1.255 0.16 1.445 0.1 1.445 0.1 1.055 0.16 1.055 0.16 1.195 0.51 1.195 0.51 1.055 0.57 1.055 0.57 1.155 0.92 1.155 0.92 1.055 0.98 1.055 0.98 1.155 1.805 1.155 ;
  END
END NOR4X4

MACRO NOR4X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X6 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5539 LAYER Metal1 ;
    ANTENNADIFFAREA 3.9397 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.535 1.37 4.475 1.37 4.475 0.98 4.125 0.98 4.125 1.21 4.065 1.21 4.065 1.15 3.65 1.15 3.65 1.21 3.59 1.21 3.59 0.92 3.65 0.92 3.65 1.09 4.065 1.09 4.065 0.92 4.26 0.92 4.26 0.64 0.33 0.64 0.33 0.35 0.39 0.35 0.39 0.58 0.74 0.58 0.74 0.35 0.8 0.35 0.8 0.58 1.15 0.58 1.15 0.35 1.21 0.35 1.21 0.58 1.615 0.58 1.615 0.35 1.675 0.35 1.675 0.58 2.025 0.58 2.025 0.35 2.085 0.35 2.085 0.58 2.545 0.58 2.545 0.35 2.605 0.35 2.605 0.58 2.955 0.58 2.955 0.35 3.015 0.35 3.015 0.58 3.365 0.58 3.365 0.35 3.425 0.35 3.425 0.58 3.87 0.58 3.87 0.35 3.93 0.35 3.93 0.58 4.28 0.58 4.28 0.35 4.34 0.35 4.34 0.73 4.32 0.73 4.32 0.92 4.475 0.92 4.475 0.9 4.535 0.9 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 0.991453 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 0.92 0.66 0.92 0.66 0.83 0.34 0.83 0.34 0.75 0.66 0.75 0.66 0.74 0.74 0.74 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 0.991453 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.835 0.84 1.575 0.84 1.575 0.895 1.435 0.895 1.435 0.84 1.39 0.84 1.39 0.76 1.835 0.76 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.24786325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.14 0.92 3.06 0.92 3.06 0.82 2.59 0.82 2.59 0.74 3.14 0.74 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 0.991453 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.125 0.82 3.965 0.82 3.965 0.895 3.835 0.895 3.835 0.82 3.7 0.82 3.7 0.74 4.125 0.74 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.125 1.65 0.125 0.9 0.185 0.9 0.185 1.65 0.535 1.65 0.535 1.25 0.595 1.25 0.595 1.65 0.945 1.65 0.945 1.25 1.005 1.25 1.005 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 4.545 0.06 4.545 0.66 4.485 0.66 4.485 0.06 4.135 0.06 4.135 0.47 4.075 0.47 4.075 0.06 3.725 0.06 3.725 0.47 3.665 0.47 3.665 0.06 3.22 0.06 3.22 0.47 3.16 0.47 3.16 0.06 2.81 0.06 2.81 0.47 2.75 0.47 2.75 0.06 2.29 0.06 2.29 0.47 2.23 0.47 2.23 0.06 1.88 0.06 1.88 0.47 1.82 0.47 1.82 0.06 1.47 0.06 1.47 0.47 1.41 0.47 1.41 0.06 1.005 0.06 1.005 0.47 0.945 0.47 0.945 0.06 0.595 0.06 0.595 0.47 0.535 0.47 0.535 0.06 0.185 0.06 0.185 0.66 0.125 0.66 0.125 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.33 1.37 3.31 1.37 3.31 1.15 2.96 1.15 2.96 1.21 2.9 1.21 2.9 0.98 2.55 0.98 2.55 1.21 2.49 1.21 2.49 0.92 2.96 0.92 2.96 1.09 3.31 1.09 3.31 0.9 3.37 0.9 3.37 1.31 3.795 1.31 3.795 1.25 3.855 1.25 3.855 1.31 4.27 1.31 4.27 1.25 4.33 1.25 ;
      POLYGON 3.165 1.37 2.23 1.37 2.23 1.055 1.88 1.055 1.88 1.21 1.82 1.21 1.82 1.055 1.415 1.055 1.415 1.21 1.355 1.21 1.355 0.995 1.82 0.995 1.82 0.94 1.88 0.94 1.88 0.995 2.23 0.995 2.23 0.9 2.29 0.9 2.29 1.31 2.695 1.31 2.695 1.25 2.755 1.25 2.755 1.31 3.105 1.31 3.105 1.25 3.165 1.25 ;
      POLYGON 2.085 1.37 1.15 1.37 1.15 1.08 0.8 1.08 0.8 1.37 0.74 1.37 0.74 1.08 0.39 1.08 0.39 1.37 0.33 1.37 0.33 0.93 0.39 0.93 0.39 1.02 1.15 1.02 1.15 0.9 1.21 0.9 1.21 1.31 1.56 1.31 1.56 1.25 1.62 1.25 1.62 1.31 2.025 1.31 2.025 1.25 2.085 1.25 ;
  END
END NOR4X6

MACRO NOR4X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4X8 0 0 ;
  SIZE 6.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.10805 LAYER Metal1 ;
    ANTENNADIFFAREA 4.929 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.935 1.345 5.875 1.345 5.875 0.875 5.54 0.875 5.54 0.92 5.525 0.92 5.525 1.185 5.46 1.185 5.46 1.055 5.115 1.055 5.115 1.185 5.055 1.185 5.055 1.055 4.705 1.055 4.705 1.185 4.645 1.185 4.645 0.995 5.3 0.995 5.3 0.815 5.46 0.815 5.46 0.79 5.49 0.79 5.49 0.53 0.335 0.53 0.335 0.515 0.26 0.515 0.26 0.455 0.38 0.455 0.38 0.47 0.67 0.47 0.67 0.455 0.79 0.455 0.79 0.47 1.08 0.47 1.08 0.455 1.2 0.455 1.2 0.47 1.49 0.47 1.49 0.455 1.61 0.455 1.61 0.47 1.95 0.47 1.95 0.455 2.07 0.455 2.07 0.47 2.36 0.47 2.36 0.455 2.48 0.455 2.48 0.47 2.77 0.47 2.77 0.455 2.89 0.455 2.89 0.47 3.18 0.47 3.18 0.455 3.3 0.455 3.3 0.47 3.59 0.47 3.59 0.455 3.71 0.455 3.71 0.47 4 0.47 4 0.455 4.12 0.455 4.12 0.47 4.41 0.47 4.41 0.455 4.53 0.455 4.53 0.47 4.82 0.47 4.82 0.455 4.94 0.455 4.94 0.47 5.23 0.47 5.23 0.455 5.35 0.455 5.35 0.47 5.67 0.47 5.67 0.41 5.73 0.41 5.73 0.53 5.55 0.53 5.55 0.815 5.935 0.815 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.081081 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.03 0.83 0.94 0.83 0.94 0.92 0.86 0.92 0.86 0.83 0.4 0.83 0.4 0.75 0.95 0.75 0.95 0.71 1.03 0.71 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.010296 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.545 0.85 2.165 0.85 2.165 0.895 2.035 0.895 2.035 0.85 1.885 0.85 1.885 0.77 2.545 0.77 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.5830115 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.34 0.92 4.26 0.92 4.26 0.83 3.32 0.83 3.32 0.77 4.225 0.77 4.225 0.71 4.285 0.71 4.285 0.77 4.34 0.77 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.15830125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.39 0.71 4.965 0.71 4.965 0.895 4.755 0.895 4.755 0.63 5.39 0.63 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 0 1.77 0 1.65 0.085 1.65 0.085 0.9 0.145 0.9 0.145 1.65 0.495 1.65 0.495 1.225 0.555 1.225 0.555 1.65 0.905 1.65 0.905 1.225 0.965 1.225 0.965 1.65 1.315 1.65 1.315 1.225 1.375 1.225 1.375 1.65 6.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 5.935 0.06 5.935 0.37 5.875 0.37 5.875 0.06 5.525 0.06 5.525 0.37 5.465 0.37 5.465 0.06 5.115 0.06 5.115 0.37 5.055 0.37 5.055 0.06 4.705 0.06 4.705 0.37 4.645 0.37 4.645 0.06 4.295 0.06 4.295 0.37 4.235 0.37 4.235 0.06 3.885 0.06 3.885 0.37 3.825 0.37 3.825 0.06 3.475 0.06 3.475 0.37 3.415 0.37 3.415 0.06 3.065 0.06 3.065 0.37 3.005 0.37 3.005 0.06 2.655 0.06 2.655 0.37 2.595 0.37 2.595 0.06 2.245 0.06 2.245 0.37 2.185 0.37 2.185 0.06 1.835 0.06 1.835 0.37 1.775 0.37 1.775 0.06 1.375 0.06 1.375 0.37 1.315 0.37 1.315 0.06 0.965 0.06 0.965 0.37 0.905 0.37 0.905 0.06 0.555 0.06 0.555 0.37 0.495 0.37 0.495 0.06 0.145 0.06 0.145 0.37 0.085 0.37 0.085 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.73 1.345 4.44 1.345 4.44 1.125 4.09 1.125 4.09 1.185 4.03 1.185 4.03 0.99 3.68 0.99 3.68 1.185 3.62 1.185 3.62 0.99 3.27 0.99 3.27 1.185 3.21 1.185 3.21 0.93 4.09 0.93 4.09 1.065 4.44 1.065 4.44 0.9 4.5 0.9 4.5 1.285 4.85 1.285 4.85 1.225 4.91 1.225 4.91 1.285 5.26 1.285 5.26 1.225 5.32 1.225 5.32 1.285 5.67 1.285 5.67 1.225 5.73 1.225 ;
      POLYGON 4.295 1.345 3.005 1.345 3.005 1.055 2.655 1.055 2.655 1.185 2.595 1.185 2.595 1.055 2.245 1.055 2.245 1.185 2.185 1.185 2.185 1.055 1.835 1.055 1.835 1.185 1.775 1.185 1.775 0.995 3.065 0.995 3.065 1.285 3.415 1.285 3.415 1.225 3.475 1.225 3.475 1.285 3.825 1.285 3.825 1.225 3.885 1.225 3.885 1.285 4.235 1.285 4.235 1.225 4.295 1.225 ;
      POLYGON 2.86 1.345 1.52 1.345 1.52 0.96 1.17 0.96 1.17 1.345 1.11 1.345 1.11 1.125 0.76 1.125 0.76 1.345 0.7 1.345 0.7 0.99 0.35 0.99 0.35 1.345 0.29 1.345 0.29 0.93 0.76 0.93 0.76 1.065 1.11 1.065 1.11 0.9 1.58 0.9 1.58 1.285 1.98 1.285 1.98 1.225 2.04 1.225 2.04 1.285 2.39 1.285 2.39 1.225 2.45 1.225 2.45 1.285 2.8 1.285 2.8 1.225 2.86 1.225 ;
  END
END NOR4X8

MACRO NOR4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3858 LAYER Metal1 ;
    ANTENNADIFFAREA 0.58715 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.11 1.04 1.11 1.04 0.98 1.08 0.98 1.08 0.545 0.35 0.545 0.35 0.29 0.41 0.29 0.41 0.485 0.79 0.485 0.79 0.29 0.85 0.29 0.85 0.485 1.14 0.485 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.36 0.895 0.03 0.895 0.03 0.815 0.125 0.815 0.125 0.645 0.36 0.645 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.73 0.54 1.23 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.645 0.74 1.145 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.98 0.73 0.94 0.73 0.94 1.11 0.86 1.11 0.86 0.65 0.98 0.65 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.145 1.65 0.145 0.995 0.205 0.995 0.205 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 1.09 0.06 1.09 0.385 1.03 0.385 1.03 0.06 0.615 0.06 0.615 0.385 0.555 0.385 0.555 0.06 0.205 0.06 0.205 0.385 0.145 0.385 0.145 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
END NOR4XL

MACRO OA21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.566 LAYER Metal1 ;
    ANTENNADIFFAREA 0.71465 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.35042725 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 145.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 0.55 1.11 0.55 1.11 0.705 0.98 0.705 0.98 1.455 0.92 1.455 0.92 0.625 1.05 0.625 1.05 0.4 1.14 0.4 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.425926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.56 0.155 0.92 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.611111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.39 1.11 0.235 1.11 0.235 0.98 0.295 0.98 0.295 0.8 0.39 0.8 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.55 0.62 0.73 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.16 0.13 1.16 0.13 1.65 0.715 1.65 0.715 1.065 0.775 1.065 0.775 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.875 0.06 0.875 0.29 0.815 0.29 0.815 0.06 0.365 0.06 0.365 0.2 0.305 0.2 0.305 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.8 0.965 0.54 0.965 0.54 1.185 0.48 1.185 0.48 0.905 0.685 0.905 0.685 0.395 0.745 0.395 0.745 0.845 0.8 0.845 ;
      RECT 0.04 0.37 0.56 0.46 ;
  END
END OA21X1

MACRO OA21X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7488 LAYER Metal1 ;
    ANTENNADIFFAREA 0.985225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.8 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 93.5384615 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.495 0.63 1.34 0.63 1.34 0.73 1.26 0.73 1.26 1.455 1.2 1.455 1.2 0.67 1.26 0.67 1.26 0.6 1.28 0.6 1.28 0.57 1.495 0.57 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.56 0.34 1.06 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.705 0.865 0.54 0.865 0.54 0.925 0.46 0.925 0.46 0.785 0.625 0.785 0.625 0.59 0.705 0.59 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.22 0.94 0.72 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.3 1.65 0.3 1.16 0.36 1.16 0.36 1.65 0.995 1.65 0.995 1.125 1.055 1.125 1.055 1.65 1.405 1.65 1.405 1.065 1.465 1.065 1.465 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.67 0.06 1.67 0.52 1.61 0.52 1.61 0.06 1.23 0.06 1.23 0.2 1.17 0.2 1.17 0.06 0.595 0.06 0.595 0.2 0.535 0.2 0.535 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.1 1.025 0.8 1.025 0.8 1.185 0.74 1.185 0.74 0.965 1.04 0.965 1.04 0.395 1.1 0.395 ;
      POLYGON 0.76 0.49 0.68 0.49 0.68 0.46 0.27 0.46 0.27 0.38 0.68 0.38 0.68 0.37 0.76 0.37 ;
  END
END OA21X2

MACRO OA21X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21X4 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.07085 LAYER Metal1 ;
    ANTENNADIFFAREA 1.415 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.152564 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 68.5384615 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 1 1.67 1 1.67 1.35 1.61 1.35 1.61 1 1.26 1 1.26 1.35 1.2 1.35 1.2 0.94 1.755 0.94 1.755 0.68 1.3 0.68 1.3 0.54 1.36 0.54 1.36 0.62 1.71 0.62 1.71 0.54 1.77 0.54 1.77 0.62 1.815 0.62 1.815 0.79 1.94 0.79 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.63 0.14 1.13 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.605 0.895 0.435 0.895 0.435 0.71 0.29 0.71 0.29 0.63 0.605 0.63 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 0.97 0.86 0.97 0.86 0.87 0.72 0.87 0.72 0.61 0.8 0.61 0.8 0.79 0.94 0.79 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.28 1.65 0.28 1.23 0.34 1.23 0.34 1.65 0.795 1.65 0.795 1.23 0.855 1.23 0.855 1.65 1.405 1.65 1.405 1.1 1.465 1.1 1.465 1.65 1.815 1.65 1.815 1.1 1.875 1.1 1.875 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 1.975 0.06 1.975 0.52 1.915 0.52 1.915 0.06 1.565 0.06 1.565 0.52 1.505 0.52 1.505 0.06 1.125 0.06 1.125 0.2 1.065 0.2 1.065 0.06 0.445 0.06 0.445 0.35 0.385 0.35 0.385 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.655 0.84 1.1 0.84 1.1 1.13 0.65 1.13 0.65 1.35 0.59 1.35 0.59 1.07 1.04 1.07 1.04 0.51 0.795 0.51 0.795 0.37 0.855 0.37 0.855 0.45 1.1 0.45 1.1 0.78 1.655 0.78 ;
      POLYGON 0.65 0.53 0.18 0.53 0.18 0.37 0.26 0.37 0.26 0.45 0.57 0.45 0.57 0.37 0.65 0.37 ;
  END
END OA21X4

MACRO OA21XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA21XL 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6366 LAYER Metal1 ;
    ANTENNADIFFAREA 0.75485 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 39.29629625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 272.4074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.38 0.65 1.34 0.65 1.34 0.73 1.13 0.73 1.13 1.185 1.05 1.185 1.05 0.65 1.26 0.65 1.26 0.57 1.38 0.57 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.56 0.34 1.06 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.22 0.74 0.72 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.185 1.65 0.185 1.16 0.245 1.16 0.245 1.65 0.845 1.65 0.845 1.16 0.905 1.16 0.905 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.185 0.06 1.185 0.2 1.125 0.2 1.125 0.06 0.395 0.06 0.395 0.2 0.335 0.2 0.335 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.95 0.845 0.9 0.845 0.9 0.88 0.7 0.88 0.7 1.185 0.64 1.185 0.64 0.82 0.84 0.82 0.84 0.395 0.9 0.395 0.9 0.725 0.95 0.725 ;
      POLYGON 0.56 0.49 0.48 0.49 0.48 0.46 0.07 0.46 0.07 0.38 0.48 0.38 0.48 0.37 0.56 0.37 ;
  END
END OA21XL

MACRO OA22X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5751 LAYER Metal1 ;
    ANTENNADIFFAREA 0.8323 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.6615385 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 157.3846155 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.73 1.305 0.73 1.305 1.33 1.245 1.33 1.245 0.37 1.305 0.37 1.305 0.41 1.34 0.41 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.4814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.805 0.87 0.94 1.085 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.79 0.39 1.015 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.83333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.2 0.775 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.4814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.87 0.57 1.11 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.21 0.13 1.21 0.13 1.65 1.04 1.65 1.04 1.21 1.1 1.21 1.1 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 1.14 0.06 1.14 0.2 1.08 0.2 1.08 0.06 0.365 0.06 0.365 0.2 0.305 0.2 0.305 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.18 0.77 0.735 0.77 0.735 1.3 0.44 1.3 0.44 1.24 0.675 1.24 0.675 0.445 0.735 0.445 0.735 0.71 1.18 0.71 ;
      POLYGON 0.94 0.54 0.88 0.54 0.88 0.345 0.53 0.345 0.53 0.54 0.47 0.54 0.47 0.51 0.04 0.51 0.04 0.45 0.47 0.45 0.47 0.285 0.94 0.285 ;
  END
END OA22X1

MACRO OA22X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8286 LAYER Metal1 ;
    ANTENNADIFFAREA 1.085025 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.1641025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 109.4358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.615 0.63 1.54 0.63 1.54 0.73 1.5 0.73 1.5 1.395 1.44 1.395 1.44 0.67 1.46 0.67 1.46 0.57 1.615 0.57 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 1.11 1.26 1.11 1.26 1.06 1.08 1.06 1.08 1.17 1 1.17 1 0.98 1.34 0.98 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.675 0.54 1.175 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.675 0.34 1.175 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.675 0.74 1.175 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.205 1.65 0.205 1.275 0.265 1.275 0.265 1.65 1.125 1.65 1.125 1.275 1.185 1.275 1.185 1.65 1.645 1.65 1.645 1.005 1.705 1.005 1.705 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.79 0.06 1.79 0.52 1.73 0.52 1.73 0.06 1.35 0.06 1.35 0.2 1.29 0.2 1.29 0.06 0.46 0.06 0.46 0.415 0.4 0.415 0.4 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.34 0.88 0.9 0.88 0.9 1.335 0.575 1.335 0.575 1.275 0.84 1.275 0.84 0.32 0.9 0.32 0.9 0.82 1.34 0.82 ;
      POLYGON 1.19 0.415 1.13 0.415 1.13 0.22 0.665 0.22 0.665 0.575 0.225 0.575 0.225 0.41 0.165 0.41 0.165 0.35 0.285 0.35 0.285 0.515 0.605 0.515 0.605 0.16 1.19 0.16 ;
  END
END OA22X2

MACRO OA22X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22X4 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.142425 LAYER Metal1 ;
    ANTENNADIFFAREA 1.5029 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.76431625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 74.4102565 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.14 1.11 1.71 1.11 1.71 1.44 1.65 1.44 1.65 1.11 1.3 1.11 1.3 1.44 1.24 1.44 1.24 1.05 1.945 1.05 1.945 0.52 1.56 0.52 1.56 0.5 1.49 0.5 1.49 0.44 1.61 0.44 1.61 0.46 1.945 0.46 1.945 0.41 2.005 0.41 2.005 0.98 2.14 0.98 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.22 1.06 1.22 1.06 1.06 1 1.06 1 0.78 1.08 0.78 1.08 0.98 1.14 0.98 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 1.2 0.46 1.2 0.46 0.88 0.48 0.88 0.48 0.72 0.56 0.72 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.72 0.34 1.22 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.72 0.74 1.22 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 1.77 0 1.77 0 1.65 0.265 1.65 0.265 1.32 0.325 1.32 0.325 1.65 1.035 1.65 1.035 1.32 1.095 1.32 1.095 1.65 1.445 1.65 1.445 1.21 1.505 1.21 1.505 1.65 1.855 1.65 1.855 1.21 1.915 1.21 1.915 1.65 2.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 0.06 2.21 0.06 2.21 0.39 2.15 0.39 2.15 0.06 1.77 0.06 1.77 0.3 1.83 0.3 1.83 0.36 1.71 0.36 1.71 0.06 1.375 0.06 1.375 0.39 1.315 0.39 1.315 0.06 0.485 0.06 0.485 0.46 0.425 0.46 0.425 0.06 0 0.06 0 -0.06 2.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.845 0.695 1.725 0.695 1.725 0.68 0.9 0.68 0.9 1.38 0.69 1.38 0.69 1.44 0.63 1.44 0.63 1.32 0.84 1.32 0.84 0.4 0.9 0.4 0.9 0.62 1.77 0.62 1.77 0.635 1.845 0.635 ;
      POLYGON 1.105 0.46 1.045 0.46 1.045 0.3 0.69 0.3 0.69 0.62 0.22 0.62 0.22 0.48 0.28 0.48 0.28 0.56 0.63 0.56 0.63 0.24 1.105 0.24 ;
  END
END OA22X4

MACRO OA22XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OA22XL 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6717 LAYER Metal1 ;
    ANTENNADIFFAREA 0.865275 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 41.462963 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 320.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.655 1.42 1.54 1.42 1.54 1.49 1.3 1.49 1.3 1.39 1.46 1.39 1.46 1.36 1.595 1.36 1.595 0.425 1.655 0.425 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.76 1.14 1.26 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 1.08 0.48 1.08 0.48 0.73 0.46 0.73 0.46 0.6 0.56 0.6 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 1.1 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.06 0.74 1.06 0.74 1.11 0.66 1.11 0.66 0.98 0.72 0.98 0.72 0.67 0.8 0.67 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.23 1.65 0.23 1.36 0.29 1.36 0.29 1.65 1.125 1.65 1.125 1.36 1.185 1.36 1.185 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.42 0.06 1.42 0.2 1.36 0.2 1.36 0.06 0.525 0.06 0.525 0.2 0.465 0.2 0.465 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.355 0.66 0.96 0.66 0.96 1.27 0.755 1.27 0.755 1.355 0.635 1.355 0.635 1.295 0.695 1.295 0.695 1.21 0.9 1.21 0.9 0.38 0.96 0.38 0.96 0.6 1.355 0.6 ;
      POLYGON 1.26 0.5 1.2 0.5 1.2 0.28 0.69 0.28 0.69 0.5 0.63 0.5 0.63 0.47 0.2 0.47 0.2 0.41 0.63 0.41 0.63 0.22 1.26 0.22 ;
  END
END OA22XL

MACRO OAI211X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X1 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.47145 LAYER Metal1 ;
    ANTENNADIFFAREA 0.71775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.945 1.45 0.86 1.45 0.86 1.12 0.515 1.12 0.515 1.45 0.455 1.45 0.455 1.06 0.865 1.06 0.865 0.24 0.925 0.24 0.925 1.15 0.945 1.15 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.055 0.885 0.145 1.11 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.74358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.685 0.365 0.92 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.20512825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.625 0.615 0.88 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.84615375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.785 0.855 0.695 0.855 0.695 0.54 0.66 0.54 0.66 0.41 0.785 0.41 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.21 0.13 1.21 0.13 1.65 0.66 1.65 0.66 1.21 0.72 1.21 0.72 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.335 0.06 0.335 0.36 0.275 0.36 0.275 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.54 0.5 0.07 0.5 0.07 0.375 0.13 0.375 0.13 0.44 0.48 0.44 0.48 0.375 0.54 0.375 ;
  END
END OAI211X1

MACRO OAI211X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X2 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1187 LAYER Metal1 ;
    ANTENNADIFFAREA 1.54645 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.13 0.515 2.015 0.515 2.015 0.695 1.34 0.695 1.34 1.06 1.81 1.06 1.81 1.345 1.75 1.345 1.75 1.12 1.4 1.12 1.4 1.345 1.34 1.345 1.34 1.12 0.7 1.12 0.7 1.345 0.64 1.345 0.64 1.06 1.26 1.06 1.26 0.98 1.28 0.98 1.28 0.635 1.955 0.635 1.955 0.455 2.13 0.455 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.745 0.895 0.54 0.895 0.54 1.11 0.46 1.11 0.46 0.815 0.745 0.815 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.12820525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.975 0.715 0.36 0.715 0.36 0.88 0.34 0.88 0.34 0.92 0.26 0.92 0.26 0.79 0.28 0.79 0.28 0.635 0.975 0.635 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.44 0.795 1.855 0.96 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.34 0.97 2.26 0.97 2.26 0.895 2.115 0.895 2.115 0.615 2.195 0.615 2.195 0.79 2.34 0.79 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 1.77 0 1.77 0 1.65 0.3 1.65 0.3 1.02 0.36 1.02 0.36 1.65 0.95 1.65 0.95 1.225 1.01 1.225 1.01 1.65 1.545 1.65 1.545 1.225 1.605 1.225 1.605 1.65 1.955 1.65 1.955 0.955 2.015 0.955 2.015 1.65 2.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 0.06 1.055 0.06 1.055 0.315 1.115 0.315 1.115 0.375 0.995 0.375 0.995 0.06 0.645 0.06 0.645 0.315 0.705 0.315 0.705 0.375 0.585 0.375 0.585 0.06 0.23 0.06 0.23 0.405 0.17 0.405 0.17 0.06 0 0.06 0 -0.06 2.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.305 0.415 2.245 0.415 2.245 0.355 1.855 0.355 1.855 0.415 1.795 0.415 1.795 0.355 1.46 0.355 1.46 0.375 1.34 0.375 1.34 0.315 1.41 0.315 1.41 0.295 2.305 0.295 ;
      POLYGON 1.68 0.515 1.61 0.515 1.61 0.535 0.41 0.535 0.41 0.415 0.47 0.415 0.47 0.475 0.82 0.475 0.82 0.415 0.88 0.415 0.88 0.475 1.56 0.475 1.56 0.455 1.68 0.455 ;
  END
END OAI211X2

MACRO OAI211X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211X4 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9092 LAYER Metal1 ;
    ANTENNADIFFAREA 2.6813 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.485 0.585 2.855 0.585 2.855 0.715 2 0.715 2 1.005 2.165 1.005 2.165 1.025 3.28 1.025 3.28 1.345 3.22 1.345 3.22 1.085 2.87 1.085 2.87 1.345 2.81 1.345 2.81 1.085 2.46 1.085 2.46 1.345 2.4 1.345 2.4 1.085 2.05 1.085 2.05 1.345 1.99 1.345 1.99 1.065 1.42 1.065 1.42 1.345 1.36 1.345 1.36 1.065 0.76 1.065 0.76 1.345 0.7 1.345 0.7 1.005 1.94 1.005 1.94 0.655 2.795 0.655 2.795 0.525 3.015 0.525 3.015 0.445 3.075 0.445 3.075 0.525 3.425 0.525 3.425 0.445 3.485 0.445 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.17948725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.605 0.815 1.375 0.895 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.4358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.685 0.715 0.34 0.715 0.34 0.92 0.26 0.92 0.26 0.72 0.22 0.72 0.22 0.66 0.305 0.66 0.305 0.655 1.685 0.655 ;
    END
  END A0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.5 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.355 0.88 3.14 0.88 3.14 0.92 3.06 0.92 3.06 0.87 2.93 0.87 2.93 0.79 3.275 0.79 3.275 0.76 3.355 0.76 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.1 0.815 2.6 0.895 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 1.77 0 1.77 0 1.65 0.185 1.65 0.185 1.02 0.245 1.02 0.245 1.65 1.05 1.65 1.05 1.225 1.11 1.225 1.11 1.65 1.725 1.65 1.725 1.225 1.785 1.225 1.785 1.65 2.195 1.65 2.195 1.225 2.255 1.225 2.255 1.65 2.605 1.65 2.605 1.225 2.665 1.225 2.665 1.65 3.015 1.65 3.015 1.225 3.075 1.225 3.075 1.65 3.425 1.65 3.425 0.96 3.485 0.96 3.485 1.65 3.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 0.06 1.755 0.06 1.755 0.335 1.815 0.335 1.815 0.395 1.695 0.395 1.695 0.06 1.345 0.06 1.345 0.335 1.405 0.335 1.405 0.395 1.285 0.395 1.285 0.06 0.935 0.06 0.935 0.335 0.995 0.335 0.995 0.395 0.875 0.395 0.875 0.06 0.525 0.06 0.525 0.335 0.585 0.335 0.585 0.395 0.465 0.395 0.465 0.06 0.145 0.06 0.145 0.425 0.085 0.425 0.085 0.06 0 0.06 0 -0.06 3.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.69 0.425 3.63 0.425 3.63 0.345 3.28 0.345 3.28 0.425 3.22 0.425 3.22 0.345 2.87 0.345 2.87 0.425 2.81 0.425 2.81 0.345 2.475 0.345 2.475 0.395 2.355 0.395 2.355 0.345 2.035 0.345 2.035 0.395 1.915 0.395 1.915 0.335 1.975 0.335 1.975 0.285 3.69 0.285 ;
      POLYGON 2.695 0.535 2.625 0.535 2.625 0.555 0.29 0.555 0.29 0.435 0.35 0.435 0.35 0.495 0.7 0.495 0.7 0.435 0.76 0.435 0.76 0.495 1.11 0.495 1.11 0.435 1.17 0.435 1.17 0.495 1.52 0.495 1.52 0.435 1.58 0.435 1.58 0.495 2.135 0.495 2.135 0.475 2.255 0.475 2.255 0.495 2.575 0.495 2.575 0.475 2.695 0.475 ;
  END
END OAI211X4

MACRO OAI211XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4751 LAYER Metal1 ;
    ANTENNADIFFAREA 0.614025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.38 1.06 1.38 1.06 1.31 0.58 1.31 0.58 1.25 1.04 1.25 1.04 0.295 1.1 0.295 1.1 1.19 1.14 1.19 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.8 0.34 1.3 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.65 0.54 1.15 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.745 1.15 0.665 1.15 0.665 0.92 0.66 0.92 0.66 0.655 0.745 0.655 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 0.94 1.1 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.245 1.65 0.245 1.51 0.305 1.51 0.305 1.65 0.845 1.65 0.845 1.51 0.905 1.51 0.905 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.465 0.06 0.465 0.39 0.405 0.39 0.405 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.7 0.385 0.64 0.385 0.64 0.55 0.23 0.55 0.23 0.385 0.17 0.385 0.17 0.325 0.29 0.325 0.29 0.49 0.58 0.49 0.58 0.325 0.7 0.325 ;
  END
END OAI211XL

MACRO OAI21X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X1 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4694 LAYER Metal1 ;
    ANTENNADIFFAREA 0.6012 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.765 1.15 0.54 1.15 0.54 1.48 0.48 1.48 0.48 1.09 0.685 1.09 0.685 0.25 0.745 0.25 0.745 1.07 0.765 1.07 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5384615 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.225 0.72 0.04 0.72 0.04 0.64 0.135 0.64 0.135 0.56 0.225 0.56 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.44 0.88 0.23 0.88 0.23 0.8 0.365 0.8 0.365 0.7 0.44 0.7 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.74358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.595 1.03 0.515 1.03 0.515 1.02 0.455 1.02 0.455 0.94 0.515 0.94 0.515 0.805 0.595 0.805 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.17 1.65 0.17 1.12 0.23 1.12 0.23 1.65 0.685 1.65 0.685 1.23 0.745 1.23 0.745 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.365 0.06 0.365 0.32 0.245 0.32 0.245 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.545 0.5 0.065 0.5 0.065 0.25 0.13 0.25 0.13 0.44 0.48 0.44 0.48 0.25 0.545 0.25 ;
  END
END OAI21X1

MACRO OAI21X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7997 LAYER Metal1 ;
    ANTENNADIFFAREA 1.1002 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.385 0.66 1.3 0.66 1.3 1.2 1.255 1.2 1.255 1.48 1.195 1.48 1.195 1.2 0.705 1.2 0.705 1.48 0.645 1.48 0.645 1.14 1.24 1.14 1.24 0.92 1.06 0.92 1.06 0.79 1.14 0.79 1.14 0.86 1.24 0.86 1.24 0.6 1.325 0.6 1.325 0.54 1.385 0.54 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.7 1.04 0.54 1.04 0.54 1.3 0.46 1.3 0.46 0.96 0.7 0.96 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.76923075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 0.92 0.86 0.92 0.86 0.86 0.345 0.86 0.345 0.78 0.94 0.78 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 0.92 1.48 0.92 1.48 1.2 1.4 1.2 1.4 0.76 1.48 0.76 1.48 0.79 1.54 0.79 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.3 1.65 0.3 1.09 0.36 1.09 0.36 1.65 0.955 1.65 0.955 1.36 1.015 1.36 1.015 1.65 1.4 1.65 1.4 1.3 1.46 1.3 1.46 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 0.91 0.06 0.91 0.52 0.85 0.52 0.85 0.06 0.5 0.06 0.5 0.52 0.44 0.52 0.44 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.59 0.52 1.53 0.52 1.53 0.44 1.115 0.44 1.115 0.68 0.235 0.68 0.235 0.54 0.295 0.54 0.295 0.62 0.645 0.62 0.645 0.54 0.705 0.54 0.705 0.62 1.055 0.62 1.055 0.38 1.59 0.38 ;
  END
END OAI21X2

MACRO OAI21X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21X4 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.352875 LAYER Metal1 ;
    ANTENNADIFFAREA 1.946 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.46 0.535 2.385 0.535 2.385 0.585 1.935 0.585 1.935 1.035 2.33 1.035 2.33 1.375 2.27 1.375 2.27 1.095 1.94 1.095 1.94 1.3 1.92 1.3 1.92 1.375 1.86 1.375 1.86 1.08 1.31 1.08 1.31 1.375 1.25 1.375 1.25 1.08 0.69 1.08 0.69 1.375 0.63 1.375 0.63 1.02 1.875 1.02 1.875 0.475 2.05 0.475 2.05 0.525 2.325 0.525 2.325 0.475 2.46 0.475 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.37179475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.265 0.91 0.435 0.91 0.435 0.815 0.68 0.815 0.68 0.83 1.265 0.83 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.65384625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 0.92 1.66 0.92 1.66 0.85 1.575 0.85 1.575 0.715 0.955 0.715 0.955 0.73 0.835 0.73 0.835 0.715 0.335 0.715 0.335 0.72 0.21 0.72 0.21 0.66 0.3 0.66 0.3 0.655 1.635 0.655 1.635 0.79 1.74 0.79 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.365 0.895 2.115 0.895 2.115 0.935 2.035 0.935 2.035 0.685 2.115 0.685 2.115 0.815 2.365 0.815 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 1.77 0 1.77 0 1.65 0.175 1.65 0.175 0.985 0.235 0.985 0.235 1.65 0.94 1.65 0.94 1.255 1 1.255 1 1.65 1.64 1.65 1.64 1.255 1.7 1.255 1.7 1.65 2.065 1.65 2.065 1.255 2.125 1.255 2.125 1.65 2.475 1.65 2.475 0.995 2.535 0.995 2.535 1.65 2.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 0.06 1.54 0.06 1.54 0.335 1.6 0.335 1.6 0.395 1.48 0.395 1.48 0.06 1.13 0.06 1.13 0.335 1.19 0.335 1.19 0.395 1.07 0.395 1.07 0.06 0.72 0.06 0.72 0.335 0.78 0.335 0.78 0.395 0.66 0.395 0.66 0.06 0.31 0.06 0.31 0.335 0.37 0.335 0.37 0.395 0.25 0.395 0.25 0.06 0 0.06 0 -0.06 2.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.635 0.425 2.575 0.425 2.575 0.365 2.225 0.365 2.225 0.425 2.165 0.425 2.165 0.365 1.775 0.365 1.775 0.555 0.075 0.555 0.075 0.435 0.135 0.435 0.135 0.495 0.485 0.495 0.485 0.435 0.545 0.435 0.545 0.495 0.895 0.495 0.895 0.435 0.955 0.435 0.955 0.495 1.305 0.495 1.305 0.435 1.365 0.435 1.365 0.495 1.715 0.495 1.715 0.305 2.635 0.305 ;
  END
END OAI21X4

MACRO OAI21XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21XL 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4397 LAYER Metal1 ;
    ANTENNADIFFAREA 0.47715 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 1.26 0.7 1.26 0.7 1.385 0.64 1.385 0.64 1.2 0.86 1.2 0.86 0.5 0.755 0.5 0.755 0.38 0.815 0.38 0.815 0.44 0.92 0.44 0.92 0.98 0.94 0.98 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.76 0.14 1.26 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.8 0.54 1.3 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.6 0.74 1.1 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.135 1.65 0.135 1.36 0.195 1.36 0.195 1.65 0.845 1.65 0.845 1.36 0.905 1.36 0.905 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.4 0.06 0.4 0.5 0.34 0.5 0.34 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.605 0.5 0.56 0.5 0.56 0.66 0.135 0.66 0.135 0.405 0.195 0.405 0.195 0.6 0.5 0.6 0.5 0.44 0.545 0.44 0.545 0.38 0.605 0.38 ;
  END
END OAI21XL

MACRO OAI221X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.669275 LAYER Metal1 ;
    ANTENNADIFFAREA 0.9939 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 1.3 1.18 1.3 1.18 1.49 1.095 1.49 1.095 1.15 0.66 1.15 0.66 1.48 0.6 1.48 0.6 1.09 1.215 1.09 1.215 0.54 1.275 0.54 1.275 0.975 1.34 0.975 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.025641 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.785 0.22 0.92 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.7 0.74 0.97 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.64102575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.425 1.11 0.26 1.11 0.26 0.98 0.345 0.98 0.345 0.92 0.425 0.92 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.7 0.94 0.97 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.25641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.15 0.92 1.06 0.92 1.06 0.595 1.14 0.595 1.14 0.78 1.15 0.78 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.13 1.65 0.13 1.2 0.19 1.2 0.19 1.65 0.91 1.65 0.91 1.225 0.97 1.225 0.97 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 0.49 0.06 0.49 0.25 0.37 0.25 0.37 0.06 0.18 0.06 0.18 0.25 0.04 0.25 0.04 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 0.57 0.43 1.105 0.49 ;
      RECT 0.205 0.56 0.9 0.62 ;
  END
END OAI221X1

MACRO OAI221X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X2 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2391 LAYER Metal1 ;
    ANTENNADIFFAREA 1.9733 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.54 0.92 2.5 0.92 2.5 1.215 2.4 1.215 2.4 1.405 2.34 1.405 2.34 1.215 1.74 1.215 1.74 1.275 1.68 1.275 1.68 1.215 0.72 1.215 0.72 1.275 0.66 1.275 0.66 1.155 2.44 1.155 2.44 0.475 2.5 0.475 2.5 0.79 2.54 0.79 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.12820525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.055 0.28 1.055 0.28 0.92 0.22 0.92 0.22 0.86 0.26 0.86 0.26 0.79 0.34 0.79 0.34 0.995 0.94 0.995 0.94 0.845 1 0.845 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.923077 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.14 1.055 1.4 1.055 1.4 0.845 1.46 0.845 1.46 0.995 2.06 0.995 2.06 0.79 2.14 0.79 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.84 0.895 0.635 0.895 0.635 0.795 0.44 0.795 0.44 0.715 0.715 0.715 0.715 0.815 0.84 0.815 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.96 0.795 1.765 0.795 1.765 0.895 1.56 0.895 1.56 0.815 1.685 0.815 1.685 0.715 1.96 0.715 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.555 2.34 1.055 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 1.77 0 1.77 0 1.65 0.35 1.65 0.35 1.285 0.41 1.285 0.41 1.65 0.985 1.65 0.985 1.315 1.105 1.315 1.105 1.375 1.045 1.375 1.045 1.65 2.105 1.65 2.105 1.315 2.225 1.315 2.225 1.375 2.165 1.375 2.165 1.65 2.6 1.65 2.6 1.02 2.66 1.02 2.66 1.65 2.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 0.06 1.13 0.06 1.13 0.455 1.07 0.455 1.07 0.06 0.72 0.06 0.72 0.455 0.66 0.455 0.66 0.06 0.17 0.06 0.17 0.455 0.11 0.455 0.11 0.06 0 0.06 0 -0.06 2.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.705 0.455 2.645 0.455 2.645 0.375 2.25 0.375 2.25 0.455 2.19 0.455 2.19 0.375 1.74 0.375 1.74 0.455 1.68 0.455 1.68 0.375 1.33 0.375 1.33 0.455 1.27 0.455 1.27 0.315 2.705 0.315 ;
      POLYGON 1.975 0.565 1.9 0.565 1.9 0.615 0.455 0.615 0.455 0.475 0.515 0.475 0.515 0.555 0.865 0.555 0.865 0.475 0.925 0.475 0.925 0.555 1.475 0.555 1.475 0.475 1.535 0.475 1.535 0.555 1.84 0.555 1.84 0.505 1.975 0.505 ;
  END
END OAI221X2

MACRO OAI221X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221X4 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.1549 LAYER Metal1 ;
    ANTENNADIFFAREA 3.252 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.34 0.92 4.3 0.92 4.3 1.13 4.185 1.13 4.185 1.46 4.125 1.46 4.125 1.27 3.775 1.27 3.775 1.46 3.715 1.46 3.715 1.27 3.105 1.27 3.105 1.33 3.045 1.33 3.045 1.27 2.485 1.27 2.485 1.33 2.425 1.33 2.425 1.27 1.51 1.27 1.51 1.33 1.45 1.33 1.45 1.27 0.63 1.27 0.63 1.33 0.57 1.33 0.57 1.21 3.715 1.21 3.715 1.07 3.775 1.07 3.775 1.21 4.125 1.21 4.125 1.07 4.24 1.07 4.24 0.675 3.805 0.675 3.805 0.535 3.865 0.535 3.865 0.615 4.215 0.615 4.215 0.535 4.3 0.535 4.3 0.79 4.34 0.79 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.9871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.755 1.055 0.28 1.055 0.28 0.92 0.22 0.92 0.22 0.86 0.26 0.86 0.26 0.79 0.34 0.79 0.34 0.995 1.01 0.995 1.01 0.935 1.07 0.935 1.07 0.995 1.695 0.995 1.695 0.91 1.755 0.91 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.9615385 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.54 1.11 2.09 1.11 2.09 0.875 2.15 0.875 2.15 1.05 2.77 1.05 2.77 0.94 2.89 0.94 2.89 1.05 3.46 1.05 3.46 0.91 3.54 0.91 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.5128205 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.475 0.835 0.765 0.835 0.765 0.895 0.615 0.895 0.615 0.775 1.475 0.775 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.0897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.165 0.895 3.035 0.895 3.035 0.835 2.47 0.835 2.47 0.775 3.12 0.775 3.12 0.815 3.165 0.815 ;
    END
  END B1
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.64 0.815 4.14 0.895 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.77 0 1.77 0 1.65 0.26 1.65 0.26 1.34 0.32 1.34 0.32 1.65 0.85 1.65 0.85 1.37 0.97 1.37 0.97 1.43 0.91 1.43 0.91 1.65 1.73 1.65 1.73 1.37 1.85 1.37 1.85 1.43 1.79 1.43 1.79 1.65 2.705 1.65 2.705 1.37 2.825 1.37 2.825 1.43 2.765 1.43 2.765 1.65 3.48 1.65 3.48 1.37 3.6 1.37 3.6 1.43 3.54 1.43 3.54 1.65 3.89 1.65 3.89 1.37 4.01 1.37 4.01 1.43 3.95 1.43 3.95 1.65 4.4 1.65 4.4 1.07 4.46 1.07 4.46 1.65 4.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 0.06 1.82 0.06 1.82 0.515 1.76 0.515 1.76 0.06 1.41 0.06 1.41 0.515 1.35 0.515 1.35 0.06 1 0.06 1 0.515 0.94 0.515 0.94 0.06 0.59 0.06 0.59 0.515 0.53 0.515 0.53 0.06 0.17 0.06 0.17 0.515 0.11 0.515 0.11 0.06 0 0.06 0 -0.06 4.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.48 0.515 4.42 0.515 4.42 0.435 4.07 0.435 4.07 0.515 4.01 0.515 4.01 0.435 3.66 0.435 3.66 0.515 3.6 0.515 3.6 0.435 3.25 0.435 3.25 0.515 3.19 0.515 3.19 0.435 2.84 0.435 2.84 0.515 2.78 0.515 2.78 0.435 2.43 0.435 2.43 0.515 2.37 0.515 2.37 0.435 2.02 0.435 2.02 0.515 1.96 0.515 1.96 0.375 4.48 0.375 ;
      POLYGON 3.485 0.625 3.41 0.625 3.41 0.675 0.325 0.675 0.325 0.535 0.385 0.535 0.385 0.615 0.735 0.615 0.735 0.535 0.795 0.535 0.795 0.615 1.145 0.615 1.145 0.535 1.205 0.535 1.205 0.615 1.555 0.615 1.555 0.535 1.615 0.535 1.615 0.615 2.165 0.615 2.165 0.535 2.225 0.535 2.225 0.615 2.575 0.615 2.575 0.535 2.635 0.535 2.635 0.615 2.985 0.615 2.985 0.535 3.045 0.535 3.045 0.615 3.35 0.615 3.35 0.565 3.485 0.565 ;
  END
END OAI221X4

MACRO OAI221XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221XL 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.756675 LAYER Metal1 ;
    ANTENNADIFFAREA 0.91945 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 1.3 1.56 1.3 1.56 1.175 0.985 1.175 0.985 1.3 0.925 1.3 0.925 1.115 1.645 1.115 1.645 0.325 1.705 0.325 1.705 1.17 1.74 1.17 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.675 0.34 1.175 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.645 0.815 1.145 0.895 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.545 1.25 0.54 1.25 0.54 1.3 0.46 1.3 0.46 1.17 0.465 1.17 0.465 0.805 0.545 0.805 ;
    END
  END A1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.515 1.34 1.015 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.52 1.545 1.015 ;
    END
  END C0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.205 1.65 0.205 1.275 0.265 1.275 0.265 1.65 1.335 1.65 1.335 1.275 1.395 1.275 1.395 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 0.65 0.06 0.65 0.2 0.59 0.2 0.59 0.06 0.25 0.06 0.25 0.2 0.19 0.2 0.19 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.52 0.42 1.44 0.42 1.44 0.255 1 0.255 1 0.39 0.88 0.39 0.88 0.31 0.92 0.31 0.92 0.175 1.52 0.175 ;
      POLYGON 1.22 0.415 1.16 0.415 1.16 0.575 0.325 0.575 0.325 0.515 1.1 0.515 1.1 0.355 1.22 0.355 ;
  END
END OAI221XL

MACRO OAI222X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X1 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.790475 LAYER Metal1 ;
    ANTENNADIFFAREA 1.1427 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 1.49 1.4 1.49 1.4 1.47 1.34 1.47 1.34 1.17 0.68 1.17 0.68 1.47 0.62 1.47 0.62 1.11 1.445 1.11 1.445 0.51 1.235 0.51 1.235 0.37 1.295 0.37 1.295 0.45 1.505 0.45 1.505 1.165 1.54 1.165 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.655 0.585 0.755 1.02 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.6153845 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.34 1.12 0.26 1.12 0.26 1.085 0.22 1.085 0.22 0.79 0.34 0.79 ;
    END
  END A0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.5128205 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.05 0.41 1.165 0.735 ;
    END
  END C0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 1.31 0.46 1.31 0.46 1.06 0.4 1.06 0.4 0.77 0.54 0.77 ;
    END
  END A1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.076923 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.74 1.365 0.935 ;
    END
  END C1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.4615385 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.95 0.93 0.86 0.93 0.86 0.585 0.94 0.585 0.94 0.78 0.95 0.78 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.145 1.65 0.145 1.145 0.205 1.145 0.205 1.65 1.03 1.65 1.03 1.23 1.09 1.23 1.09 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 0.51 0.06 0.51 0.23 0.39 0.23 0.39 0.06 0.175 0.06 0.175 0.23 0.055 0.23 0.055 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.5 0.35 1.44 0.35 1.44 0.27 1.09 0.27 1.09 0.35 1.03 0.35 1.03 0.27 0.68 0.27 0.68 0.35 0.62 0.35 0.62 0.21 1.5 0.21 ;
      POLYGON 0.885 0.49 0.31 0.49 0.31 0.66 0.25 0.66 0.25 0.43 0.825 0.43 0.825 0.37 0.885 0.37 ;
  END
END OAI222X1

MACRO OAI222X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X2 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4924 LAYER Metal1 ;
    ANTENNADIFFAREA 2.2642 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.34 0.73 3.32 0.73 3.32 1.215 2.58 1.215 2.58 1.275 2.52 1.275 2.52 1.215 1.745 1.215 1.745 1.275 1.685 1.275 1.685 1.215 0.685 1.215 0.685 1.275 0.625 1.275 0.625 1.155 3.26 1.155 3.26 0.555 2.415 0.555 2.415 0.415 2.475 0.415 2.475 0.495 2.825 0.495 2.825 0.415 2.885 0.415 2.885 0.495 3.32 0.495 3.32 0.6 3.34 0.6 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.5384615 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 1.055 0.275 1.055 0.275 0.845 0.335 0.845 0.335 0.995 0.86 0.995 0.86 0.79 0.94 0.79 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.82051275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.14 1.055 1.46 1.055 1.46 0.895 1.42 0.895 1.42 0.835 1.46 0.835 1.46 0.79 1.54 0.79 1.54 0.995 2.08 0.995 2.08 0.845 2.14 0.845 ;
    END
  END B0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.82051275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.98 0.85 2.94 0.85 2.94 0.92 2.92 0.92 2.92 1.055 2.26 1.055 2.26 0.845 2.32 0.845 2.32 0.995 2.86 0.995 2.86 0.79 2.98 0.79 ;
    END
  END C0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.675 0.65 0.895 ;
    END
  END A1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.76 0.895 2.42 0.895 2.42 0.775 2.68 0.775 2.68 0.655 2.76 0.655 ;
    END
  END C1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.98 0.895 1.835 0.895 1.835 0.735 1.64 0.735 1.64 0.655 1.98 0.655 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 1.77 0 1.77 0 1.65 0.2 1.65 0.2 1.285 0.26 1.285 0.26 1.65 0.96 1.65 0.96 1.315 1.08 1.315 1.08 1.375 1.02 1.375 1.02 1.65 2.18 1.65 2.18 1.315 2.3 1.315 2.3 1.375 2.24 1.375 2.24 1.65 2.8 1.65 2.8 1.315 2.92 1.315 2.92 1.375 2.86 1.375 2.86 1.65 3.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 0.06 1.05 0.06 1.05 0.395 0.99 0.395 0.99 0.06 0.615 0.06 0.615 0.395 0.555 0.395 0.555 0.06 0.205 0.06 0.205 0.395 0.145 0.395 0.145 0.06 0 0.06 0 -0.06 3.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.09 0.395 3.03 0.395 3.03 0.315 2.68 0.315 2.68 0.395 2.62 0.395 2.62 0.315 2.27 0.315 2.27 0.395 2.21 0.395 2.21 0.315 1.79 0.315 1.79 0.395 1.73 0.395 1.73 0.315 1.38 0.315 1.38 0.395 1.32 0.395 1.32 0.255 3.09 0.255 ;
      POLYGON 1.995 0.555 0.35 0.555 0.35 0.415 0.41 0.415 0.41 0.495 0.76 0.495 0.76 0.415 0.82 0.415 0.82 0.495 1.525 0.495 1.525 0.415 1.585 0.415 1.585 0.495 1.935 0.495 1.935 0.415 1.995 0.415 ;
  END
END OAI222X2

MACRO OAI222X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222X4 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.460475 LAYER Metal1 ;
    ANTENNADIFFAREA 3.73675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.14 0.92 5.12 0.92 5.12 1.215 4.69 1.215 4.69 1.275 4.63 1.275 4.63 1.215 4.065 1.215 4.065 1.275 4.005 1.275 4.005 1.215 3.28 1.215 3.28 1.275 3.22 1.275 3.22 1.215 2.425 1.215 2.425 1.275 2.365 1.275 2.365 1.215 1.505 1.215 1.505 1.275 1.445 1.275 1.445 1.215 0.835 1.215 0.835 1.275 0.775 1.275 0.775 1.155 5.06 1.155 5.06 0.675 3.835 0.675 3.835 0.535 3.895 0.535 3.895 0.615 4.245 0.615 4.245 0.535 4.305 0.535 4.305 0.615 4.655 0.615 4.655 0.535 4.715 0.535 4.715 0.615 5.065 0.615 5.065 0.535 5.125 0.535 5.125 0.79 5.14 0.79 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 1.055 0.305 1.055 0.305 0.935 0.365 0.935 0.365 0.995 1.065 0.995 1.065 0.935 1.185 0.935 1.185 0.995 1.66 0.995 1.66 0.79 1.74 0.79 ;
    END
  END A0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.15384625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.925 1.055 3.86 1.055 3.86 0.895 3.73 0.895 3.73 0.835 3.86 0.835 3.86 0.79 3.94 0.79 3.94 0.995 4.35 0.995 4.35 0.935 4.47 0.935 4.47 0.995 4.865 0.995 4.865 0.895 4.925 0.895 ;
    END
  END C0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.82051275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.54 0.92 3.52 0.92 3.52 1.055 2.085 1.055 2.085 0.895 2.145 0.895 2.145 0.995 2.685 0.995 2.685 0.935 2.805 0.935 2.805 0.995 3.46 0.995 3.46 0.79 3.54 0.79 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.35897425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.47 0.835 0.965 0.835 0.965 0.895 0.835 0.895 0.835 0.835 0.67 0.835 0.67 0.775 1.47 0.775 ;
    END
  END A1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.16666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.765 0.895 4.635 0.895 4.635 0.835 4.04 0.835 4.04 0.775 4.765 0.775 ;
    END
  END C1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.21794875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.18 0.835 2.585 0.835 2.585 0.895 2.435 0.895 2.435 0.775 3.18 0.775 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 1.77 0 1.77 0 1.65 0.465 1.65 0.465 1.335 0.525 1.335 0.525 1.65 1.105 1.65 1.105 1.365 1.225 1.365 1.225 1.425 1.165 1.425 1.165 1.65 1.725 1.65 1.725 1.365 1.845 1.365 1.845 1.425 1.785 1.425 1.785 1.65 2.825 1.65 2.825 1.365 2.945 1.365 2.945 1.425 2.885 1.425 2.885 1.65 3.525 1.65 3.525 1.365 3.645 1.365 3.645 1.425 3.585 1.425 3.585 1.65 4.285 1.65 4.285 1.365 4.405 1.365 4.405 1.425 4.345 1.425 4.345 1.65 4.91 1.65 4.91 1.365 5.03 1.365 5.03 1.425 4.97 1.425 4.97 1.65 5.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 0.06 1.815 0.06 1.815 0.515 1.755 0.515 1.755 0.06 1.405 0.06 1.405 0.515 1.345 0.515 1.345 0.06 0.995 0.06 0.995 0.515 0.935 0.515 0.935 0.06 0.585 0.06 0.585 0.515 0.525 0.515 0.525 0.06 0.175 0.06 0.175 0.515 0.115 0.515 0.115 0.06 0 0.06 0 -0.06 5.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.33 0.515 5.27 0.515 5.27 0.435 4.92 0.435 4.92 0.515 4.86 0.515 4.86 0.435 4.51 0.435 4.51 0.515 4.45 0.515 4.45 0.435 4.1 0.435 4.1 0.515 4.04 0.515 4.04 0.435 3.69 0.435 3.69 0.515 3.63 0.515 3.63 0.435 3.28 0.435 3.28 0.515 3.22 0.515 3.22 0.435 2.84 0.435 2.84 0.515 2.78 0.515 2.78 0.435 2.425 0.435 2.425 0.515 2.365 0.515 2.365 0.435 2.015 0.435 2.015 0.515 1.955 0.515 1.955 0.375 5.33 0.375 ;
      POLYGON 3.485 0.675 0.32 0.675 0.32 0.535 0.38 0.535 0.38 0.615 0.73 0.615 0.73 0.535 0.79 0.535 0.79 0.615 1.14 0.615 1.14 0.535 1.2 0.535 1.2 0.615 1.55 0.615 1.55 0.535 1.61 0.535 1.61 0.615 2.16 0.615 2.16 0.535 2.22 0.535 2.22 0.615 2.57 0.615 2.57 0.535 2.63 0.535 2.63 0.615 2.985 0.615 2.985 0.535 3.045 0.535 3.045 0.615 3.425 0.615 3.425 0.535 3.485 0.535 ;
  END
END OAI222X4

MACRO OAI222XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222XL 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.753275 LAYER Metal1 ;
    ANTENNADIFFAREA 0.840525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 1.315 1.345 1.315 1.345 1.23 0.66 1.23 0.66 1.31 0.6 1.31 0.6 1.165 1.45 1.165 1.45 0.68 1.245 0.68 1.245 0.465 1.305 0.465 1.305 0.62 1.51 0.62 1.51 1.165 1.54 1.165 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.24074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.76 0.76 1.105 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.99 0.22 1.15 ;
    END
  END A0
  PIN C0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.24074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.16 0.885 1.14 0.885 1.14 1.085 1.06 1.085 1.06 0.74 1.16 0.74 ;
    END
  END C0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.345 0.765 0.545 0.92 ;
    END
  END A1
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.0555555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.37 0.88 1.34 0.88 1.34 1.085 1.26 1.085 1.26 0.76 1.37 0.76 ;
    END
  END C1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.425926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.97 0.88 0.94 0.88 0.94 1.105 0.86 1.105 0.86 0.76 0.97 0.76 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.13 1.65 0.13 1.285 0.19 1.285 0.19 1.65 0.955 1.65 0.955 1.315 1.075 1.315 1.075 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 0.53 0.06 0.53 0.2 0.47 0.2 0.47 0.06 0.16 0.06 0.16 0.2 0.1 0.2 0.1 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.54 0.53 1.42 0.53 1.42 0.38 1.07 0.38 1.07 0.68 0.645 0.68 0.645 0.53 0.57 0.53 0.57 0.47 0.705 0.47 0.705 0.62 1.01 0.62 1.01 0.32 1.48 0.32 1.48 0.47 1.54 0.47 ;
      POLYGON 0.865 0.56 0.805 0.56 0.805 0.38 0.295 0.38 0.295 0.56 0.235 0.56 0.235 0.32 0.865 0.32 ;
  END
END OAI222XL

MACRO OAI22X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4731 LAYER Metal1 ;
    ANTENNADIFFAREA 0.8089 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.77 0.64 0.7 0.64 0.7 0.81 0.545 0.81 0.545 1.46 0.465 1.46 0.465 0.75 0.64 0.75 0.64 0.58 0.71 0.58 0.71 0.4 0.77 0.4 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.5641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.285 0.72 0.365 1.085 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.145 1.085 0.065 1.085 0.065 0.84 0.055 0.84 0.055 0.72 0.145 0.72 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.4102565 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.865 0.74 0.945 1.09 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.30769225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.645 0.91 0.725 1.25 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.21 0.13 1.21 0.13 1.65 0.89 1.65 0.89 1.2 0.95 1.2 0.95 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.305 0.06 0.305 0.43 0.365 0.43 0.365 0.49 0.245 0.49 0.245 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.975 0.64 0.915 0.64 0.915 0.34 0.54 0.34 0.54 0.65 0.07 0.65 0.07 0.4 0.13 0.4 0.13 0.59 0.48 0.59 0.48 0.28 0.975 0.28 ;
  END
END OAI22X1

MACRO OAI22X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.90935 LAYER Metal1 ;
    ANTENNADIFFAREA 1.3536 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.655 0.505 1.58 0.505 1.58 0.555 1.16 0.555 1.16 0.685 0.995 0.685 0.995 1.025 1.465 1.025 1.465 1.355 1.405 1.355 1.405 1.085 0.7 1.085 0.7 1.355 0.64 1.355 0.64 1.025 0.835 1.025 0.835 1.005 0.935 1.005 0.935 0.625 1.1 0.625 1.1 0.445 1.245 0.445 1.245 0.495 1.52 0.495 1.52 0.445 1.655 0.445 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.655 0.885 0.34 0.885 0.34 1.11 0.26 1.11 0.26 0.805 0.655 0.805 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 1.115 1.66 1.115 1.66 0.915 1.44 0.915 1.44 0.835 1.74 0.835 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.87179475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.835 0.745 0.755 0.745 0.755 0.705 0.2 0.705 0.2 0.625 0.835 0.625 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.6153845 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.73 0.735 1.34 0.735 1.34 0.92 1.26 0.92 1.26 0.865 1.095 0.865 1.095 0.785 1.26 0.785 1.26 0.655 1.73 0.655 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.33 1.65 0.33 1.235 0.39 1.235 0.39 1.65 0.95 1.65 0.95 1.235 1.01 1.235 1.01 1.65 1.84 1.65 1.84 0.965 1.9 0.965 1.9 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 0.765 0.06 0.765 0.305 0.825 0.305 0.825 0.365 0.705 0.365 0.705 0.06 0.325 0.06 0.325 0.305 0.385 0.305 0.385 0.365 0.265 0.365 0.265 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.83 0.395 1.77 0.395 1.77 0.335 1.42 0.335 1.42 0.395 1.36 0.395 1.36 0.335 1 0.335 1 0.525 0.115 0.525 0.115 0.505 0.045 0.505 0.045 0.445 0.165 0.445 0.165 0.465 0.485 0.465 0.485 0.445 0.605 0.445 0.605 0.465 0.94 0.465 0.94 0.275 1.83 0.275 ;
  END
END OAI22X2

MACRO OAI22X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22X4 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7208 LAYER Metal1 ;
    ANTENNADIFFAREA 2.66565 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.555 0.505 3.48 0.505 3.48 0.555 1.975 0.555 1.975 1.095 3.025 1.095 3.025 0.975 3.085 0.975 3.085 1.345 3.025 1.345 3.025 1.155 2.465 1.155 2.465 1.215 2.405 1.215 2.405 1.155 2.165 1.155 2.165 1.275 2.035 1.275 2.035 1.155 1.595 1.155 1.595 1.345 1.535 1.345 1.535 1.155 0.91 1.155 0.91 1.345 0.85 1.345 0.85 0.995 0.91 0.995 0.91 1.095 1.535 1.095 1.535 0.995 1.595 0.995 1.595 1.095 1.915 1.095 1.915 0.495 2.205 0.495 2.205 0.445 2.325 0.445 2.325 0.495 2.615 0.495 2.615 0.445 2.735 0.445 2.735 0.495 3.025 0.495 3.025 0.445 3.145 0.445 3.145 0.495 3.42 0.495 3.42 0.445 3.555 0.445 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.12820525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.745 0.815 1.495 0.895 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.102564 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.18 0.875 2.765 0.875 2.765 0.895 2.44 0.895 2.44 0.815 3.18 0.815 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.397436 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.815 0.705 0.18 0.705 0.18 0.645 1.235 0.645 1.235 0.625 1.365 0.625 1.365 0.645 1.815 0.645 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.576923 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.595 0.715 2.34 0.715 2.34 0.92 2.26 0.92 2.26 0.715 2.075 0.715 2.075 0.655 3.595 0.655 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 1.77 0 1.77 0 1.65 0.54 1.65 0.54 0.955 0.6 0.955 0.6 1.65 1.13 1.65 1.13 1.255 1.25 1.255 1.25 1.315 1.19 1.315 1.19 1.65 1.865 1.65 1.865 1.375 1.985 1.375 1.985 1.435 1.925 1.435 1.925 1.65 2.685 1.65 2.685 1.255 2.805 1.255 2.805 1.315 2.745 1.315 2.745 1.65 3.335 1.65 3.335 0.955 3.395 0.955 3.395 1.65 3.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 0.06 1.745 0.06 1.745 0.16 1.805 0.16 1.805 0.22 1.685 0.22 1.685 0.06 1.275 0.06 1.275 0.16 1.335 0.16 1.335 0.22 1.215 0.22 1.215 0.06 0.805 0.06 0.805 0.16 0.865 0.16 0.865 0.22 0.745 0.22 0.745 0.06 0.335 0.06 0.335 0.16 0.395 0.16 0.395 0.22 0.275 0.22 0.275 0.06 0 0.06 0 -0.06 3.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.73 0.395 3.67 0.395 3.67 0.335 3.32 0.335 3.32 0.395 3.26 0.395 3.26 0.335 2.91 0.335 2.91 0.395 2.85 0.395 2.85 0.335 2.5 0.335 2.5 0.395 2.44 0.395 2.44 0.335 2.01 0.335 2.01 0.395 0.04 0.395 0.04 0.335 1.95 0.335 1.95 0.275 3.73 0.275 ;
  END
END OAI22X4

MACRO OAI22XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4359 LAYER Metal1 ;
    ANTENNADIFFAREA 0.610275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.795 0.51 0.695 0.51 0.695 0.7 0.54 0.7 0.54 1.235 0.48 1.235 0.48 1.11 0.46 1.11 0.46 0.98 0.48 0.98 0.48 0.64 0.635 0.64 0.635 0.45 0.735 0.45 0.735 0.39 0.795 0.39 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.37 0.92 0.34 0.92 0.34 1.05 0.26 1.05 0.26 0.79 0.29 0.79 0.29 0.58 0.37 0.58 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 1.1 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.61 0.94 1.11 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.8 0.74 1.3 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.075 1.65 0.075 1.21 0.135 1.21 0.135 1.65 0.935 1.65 0.935 1.21 0.995 1.21 0.995 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.37 0.06 0.37 0.2 0.31 0.2 0.31 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.05 0.51 0.99 0.51 0.99 0.29 0.535 0.29 0.535 0.51 0.475 0.51 0.475 0.48 0.045 0.48 0.045 0.42 0.475 0.42 0.475 0.23 1.05 0.23 ;
  END
END OAI22XL

MACRO OAI2BB1X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X1 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.444675 LAYER Metal1 ;
    ANTENNADIFFAREA 0.61765 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 15.202564 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 129.69230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.335 1.34 0.275 1.34 0.275 1.03 0.06 1.03 0.06 0.41 0.17 0.41 0.17 0.26 0.23 0.26 0.23 0.54 0.12 0.54 0.12 0.97 0.335 0.97 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.20512825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.465 0.895 0.23 0.895 0.23 0.81 0.405 0.81 0.405 0.72 0.465 0.72 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.645 1.12 0.435 1.12 0.435 0.97 0.555 0.97 0.555 0.77 0.645 0.77 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.845 0.59 0.94 0.92 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.1 0.13 1.1 0.13 1.65 0.48 1.65 0.48 1.22 0.54 1.22 0.54 1.65 0.85 1.65 0.85 1.51 0.91 1.51 0.91 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.54 0.06 0.54 0.52 0.48 0.52 0.48 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.9 0.52 0.785 0.52 0.785 1.34 0.685 1.34 0.685 1.215 0.725 1.215 0.725 0.66 0.26 0.66 0.26 0.745 0.2 0.745 0.2 0.6 0.725 0.6 0.725 0.43 0.805 0.43 0.805 0.395 0.9 0.395 ;
  END
END OAI2BB1X1

MACRO OAI2BB1X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7901 LAYER Metal1 ;
    ANTENNADIFFAREA 1.06585 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.505983 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 99.3846155 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.86 1.48 0.8 1.48 0.8 1.17 0.45 1.17 0.45 1.48 0.39 1.48 0.39 1.17 0.06 1.17 0.06 0.98 0.17 0.98 0.17 0.61 0.595 0.61 0.595 0.53 0.655 0.53 0.655 0.67 0.23 0.67 0.23 1.11 0.86 1.11 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.79487175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.92 0.85 0.54 0.85 0.54 0.92 0.46 0.92 0.46 0.85 0.33 0.85 0.33 0.77 0.92 0.77 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.375 0.85 1.085 0.85 1.085 0.705 1.02 0.705 1.02 0.625 1.165 0.625 1.165 0.77 1.375 0.77 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 1.3 1.66 1.3 1.66 1.25 1.635 1.25 1.635 0.825 1.715 0.825 1.715 1.17 1.74 1.17 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.185 1.65 0.185 1.36 0.245 1.36 0.245 1.65 0.595 1.65 0.595 1.36 0.655 1.36 0.655 1.65 1.035 1.65 1.035 1.51 1.095 1.51 1.095 1.65 1.465 1.65 1.465 1.51 1.525 1.51 1.525 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 0.965 0.06 0.965 0.51 0.905 0.51 0.905 0.06 0.345 0.06 0.345 0.51 0.285 0.51 0.285 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.595 0.62 1.535 0.62 1.535 1.01 1.36 1.01 1.36 1.21 1.3 1.21 1.3 1.01 0.64 1.01 0.64 0.95 1.475 0.95 1.475 0.56 1.595 0.56 ;
  END
END OAI2BB1X2

MACRO OAI2BB1X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1X4 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2721 LAYER Metal1 ;
    ANTENNADIFFAREA 1.7914 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.8726495 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 82.5128205 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.635 1.44 1.575 1.44 1.575 1.22 1.225 1.22 1.225 1.44 1.165 1.44 1.165 1.22 0.805 1.22 0.805 1.44 0.745 1.44 0.745 1.22 0.395 1.22 0.395 1.44 0.335 1.44 0.335 1.22 0.06 1.22 0.06 0.98 0.115 0.98 0.115 0.59 0.51 0.59 0.51 0.57 0.63 0.57 0.63 0.59 1.095 0.59 1.095 0.57 1.36 0.57 1.36 0.63 1.145 0.63 1.145 0.65 0.175 0.65 0.175 1.16 1.635 1.16 ;
    END
  END Y
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.1 0.9 1.885 0.9 1.885 0.705 1.795 0.705 1.795 0.625 1.965 0.625 1.965 0.82 2.1 0.82 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.54 1.16 2.46 1.16 2.46 1.06 2.36 1.06 2.36 0.76 2.44 0.76 2.44 0.98 2.54 0.98 ;
    END
  END A1N
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.076923 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.695 0.81 0.54 0.81 0.54 0.92 0.46 0.92 0.46 0.81 0.275 0.81 0.275 0.75 1.695 0.75 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 1.77 0 1.77 0 1.65 0.13 1.65 0.13 1.32 0.19 1.32 0.19 1.65 0.54 1.65 0.54 1.32 0.6 1.32 0.6 1.65 0.96 1.65 0.96 1.32 1.02 1.32 1.02 1.65 1.37 1.65 1.37 1.32 1.43 1.32 1.43 1.65 1.78 1.65 1.78 1.16 1.84 1.16 1.84 1.65 2.36 1.65 2.36 1.26 2.42 1.26 2.42 1.65 2.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 0.06 1.84 0.06 1.84 0.52 1.78 0.52 1.78 0.06 0.935 0.06 0.935 0.43 0.995 0.43 0.995 0.49 0.875 0.49 0.875 0.06 0.26 0.06 0.26 0.43 0.32 0.43 0.32 0.49 0.2 0.49 0.2 0.06 0 0.06 0 -0.06 2.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.26 1.06 2.215 1.06 2.215 1.44 2.155 1.44 2.155 1.06 0.7 1.06 0.7 0.97 0.64 0.97 0.64 0.91 0.76 0.91 0.76 1 1.265 1 1.265 0.91 1.385 0.91 1.385 1 2.2 1 2.2 0.54 2.26 0.54 ;
  END
END OAI2BB1X4

MACRO OAI2BB1XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB1XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5264 LAYER Metal1 ;
    ANTENNADIFFAREA 0.597775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 32.49382725 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 248.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.47 1.34 0.41 1.34 0.41 1.28 0.3 1.28 0.3 0.68 0.08 0.68 0.08 0.54 0.06 0.54 0.06 0.41 0.08 0.41 0.08 0.3 0.28 0.3 0.28 0.24 0.34 0.24 0.34 0.36 0.14 0.36 0.14 0.62 0.36 0.62 0.36 1.22 0.47 1.22 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.62 0.54 1.12 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.62 0.74 1.12 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.61 1.14 1.11 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.245 1.65 0.245 1.51 0.305 1.51 0.305 1.65 0.645 1.65 0.645 1.51 0.705 1.51 0.705 1.65 1.005 1.65 1.005 1.51 1.065 1.51 1.065 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.65 0.06 0.65 0.36 0.59 0.36 0.59 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.975 0.51 0.9 0.51 0.9 1.245 0.84 1.245 0.84 0.52 0.315 0.52 0.315 0.46 0.84 0.46 0.84 0.45 0.915 0.45 0.915 0.265 0.975 0.265 ;
  END
END OAI2BB1XL

MACRO OAI2BB2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X1 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2116 LAYER Metal1 ;
    ANTENNADIFFAREA 1.308375 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 20.711111 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 161.5384615 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.1 1.255 1.805 1.255 1.805 1.315 1.745 1.315 1.745 1.275 1.435 1.275 1.435 1.195 2.04 1.195 2.04 0.5 1.995 0.5 1.995 0.38 2.055 0.38 2.055 0.44 2.1 0.44 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.34 0.905 2.2 0.905 2.2 0.755 2.26 0.755 2.26 0.465 2.34 0.465 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.595 1.94 1.095 ;
    END
  END B1
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.915 1.105 0.625 1.105 0.625 0.815 0.71 0.815 0.71 1.005 0.915 1.005 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.525 1.105 0.445 1.105 0.445 0.895 0.235 0.895 0.235 0.815 0.525 0.815 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 1.77 0 1.77 0 1.65 0.52 1.65 0.52 1.205 0.58 1.205 0.58 1.65 1.275 1.65 1.275 0.925 1.335 0.925 1.335 1.65 2.2 1.65 2.2 1.005 2.26 1.005 2.26 1.65 2.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 0.06 1.57 0.06 1.57 0.275 1.63 0.275 1.63 0.335 1.51 0.335 1.51 0.06 0.605 0.06 0.605 0.555 0.545 0.555 0.545 0.06 0 0.06 0 -0.06 2.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.26 0.365 2.2 0.365 2.2 0.28 1.85 0.28 1.85 0.495 1.335 0.495 1.335 0.375 1.395 0.375 1.395 0.435 1.73 0.435 1.73 0.415 1.79 0.415 1.79 0.22 2.26 0.22 ;
      POLYGON 1.76 0.655 1.175 0.655 1.175 0.365 0.765 0.365 0.765 0.715 0.135 0.715 0.135 1.11 0.345 1.11 0.345 1.23 0.285 1.23 0.285 1.17 0.075 1.17 0.075 0.655 0.315 0.655 0.315 0.465 0.375 0.465 0.375 0.655 0.705 0.655 0.705 0.305 1.235 0.305 1.235 0.595 1.76 0.595 ;
      POLYGON 1.49 0.815 1.075 0.815 1.075 1.265 0.785 1.265 0.785 1.325 0.725 1.325 0.725 1.205 1.015 1.205 1.015 0.585 0.865 0.585 0.865 0.465 0.925 0.465 0.925 0.525 1.075 0.525 1.075 0.755 1.49 0.755 ;
  END
END OAI2BB2X1

MACRO OAI2BB2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X2 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5492 LAYER Metal1 ;
    ANTENNADIFFAREA 1.979875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.24102575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 101.84615375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.81 0.46 2.735 0.46 2.735 0.64 2.135 0.64 2.135 1.205 2.53 1.205 2.53 1.325 2.47 1.325 2.47 1.265 2.075 1.265 2.075 1.085 1.7 1.085 1.7 1.455 1.64 1.455 1.64 1.085 1.435 1.085 1.435 1.005 1.565 1.005 1.565 1.025 2.075 1.025 2.075 0.58 2.28 0.58 2.28 0.4 2.4 0.4 2.4 0.46 2.34 0.46 2.34 0.58 2.675 0.58 2.675 0.4 2.81 0.4 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.84 0.945 2.635 0.945 2.635 0.895 2.465 0.895 2.465 0.815 2.635 0.815 2.635 0.74 2.84 0.74 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.87179475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3 1.105 2.235 1.105 2.235 0.775 2.295 0.775 2.295 0.815 2.365 0.815 2.365 0.895 2.295 0.895 2.295 1.045 2.94 1.045 2.94 0.87 3 0.87 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.725 0.895 0.415 0.895 0.415 0.815 0.645 0.815 0.645 0.625 0.725 0.625 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.545 0.705 0.315 0.705 0.315 0.895 0.235 0.895 0.235 0.625 0.545 0.625 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 1.77 0 1.77 0 1.65 0.385 1.65 0.385 0.995 0.445 0.995 0.445 1.65 1.275 1.65 1.275 1.065 1.335 1.065 1.335 1.65 2.035 1.65 2.035 1.365 2.155 1.365 2.155 1.425 2.095 1.425 2.095 1.65 2.78 1.65 2.78 1.335 2.84 1.335 2.84 1.65 3.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 0.06 1.89 0.06 1.89 0.26 1.95 0.26 1.95 0.32 1.83 0.32 1.83 0.06 1.45 0.06 1.45 0.26 1.51 0.26 1.51 0.32 1.39 0.32 1.39 0.06 0.535 0.06 0.535 0.365 0.475 0.365 0.475 0.06 0 0.06 0 -0.06 3.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.13 0.36 3.07 0.36 3.07 0.3 2.575 0.3 2.575 0.36 2.515 0.36 2.515 0.3 2.125 0.3 2.125 0.48 1.24 0.48 1.24 0.46 1.17 0.46 1.17 0.4 1.29 0.4 1.29 0.42 1.61 0.42 1.61 0.4 1.73 0.4 1.73 0.42 2.065 0.42 2.065 0.24 3.13 0.24 ;
      POLYGON 1.975 0.81 0.885 0.81 0.885 1.02 0.825 1.02 0.825 0.395 0.885 0.395 0.885 0.75 1.975 0.75 ;
      POLYGON 1.59 0.64 0.985 0.64 0.985 0.295 0.695 0.295 0.695 0.525 0.135 0.525 0.135 0.995 0.24 0.995 0.24 1.115 0.18 1.115 0.18 1.055 0.075 1.055 0.075 0.465 0.125 0.465 0.125 0.395 0.185 0.395 0.185 0.465 0.635 0.465 0.635 0.235 1.045 0.235 1.045 0.58 1.59 0.58 ;
  END
END OAI2BB2X2

MACRO OAI2BB2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2X4 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.84275 LAYER Metal1 ;
    ANTENNADIFFAREA 3.55635 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.234 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.14850425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 93.025641 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.67 0.365 4.55 0.365 4.55 0.345 4.23 0.345 4.23 0.365 4.11 0.365 4.11 0.345 3.675 0.345 3.675 0.365 3.615 0.365 3.615 0.525 2.965 0.525 2.965 1.215 3.465 1.215 3.465 1.155 4.45 1.155 4.45 1.215 3.525 1.215 3.525 1.275 2.485 1.275 2.485 1.335 2.425 1.335 2.425 1.17 1.765 1.17 1.765 1.23 1.705 1.23 1.705 1.11 2.735 1.11 2.735 1.215 2.835 1.215 2.835 1.195 2.905 1.195 2.905 0.465 3.115 0.465 3.115 0.445 3.235 0.445 3.235 0.465 3.555 0.465 3.555 0.305 3.625 0.305 3.625 0.285 4.6 0.285 4.6 0.305 4.67 0.305 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0584 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 0.49914525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.64102575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.545 0.705 3.365 0.705 3.365 0.745 3.285 0.745 3.285 0.705 3.085 0.705 3.085 0.625 3.545 0.625 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.79487175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.685 0.895 4.535 0.895 4.535 0.905 3.365 0.905 3.365 1.085 3.125 1.085 3.125 0.905 3.065 0.905 3.065 0.845 4.475 0.845 4.475 0.835 4.685 0.835 ;
    END
  END B0
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.685 0.54 1.185 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.685 0.34 1.185 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 1.77 0 1.77 0 1.65 0.385 1.65 0.385 1.285 0.445 1.285 0.445 1.65 1.385 1.65 1.385 1.245 1.445 1.245 1.445 1.65 2.025 1.65 2.025 1.49 2.145 1.49 2.145 1.55 2.085 1.55 2.085 1.65 2.895 1.65 2.895 1.54 3.015 1.54 3.015 1.65 3.92 1.65 3.92 1.49 4.04 1.49 4.04 1.55 3.98 1.55 3.98 1.65 4.67 1.65 4.67 1.49 4.79 1.49 4.79 1.55 4.73 1.55 4.73 1.65 5 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 0.06 2.75 0.06 2.75 0.17 2.63 0.17 2.63 0.06 2.25 0.06 2.25 0.305 2.31 0.305 2.31 0.365 2.19 0.365 2.19 0.06 1.84 0.06 1.84 0.305 1.9 0.305 1.9 0.365 1.78 0.365 1.78 0.06 1.445 0.06 1.445 0.395 1.385 0.395 1.385 0.06 0.41 0.06 0.41 0.425 0.35 0.425 0.35 0.06 0 0.06 0 -0.06 5 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.845 1.375 3.685 1.375 3.685 1.44 2.795 1.44 2.795 1.495 2.265 1.495 2.265 1.39 1.545 1.39 1.545 1.145 0.83 1.145 0.83 0.715 1.005 0.715 1.005 0.445 1.125 0.445 1.125 0.505 1.065 0.505 1.065 0.715 1.27 0.715 1.27 0.765 1.59 0.765 1.59 0.415 1.65 0.415 1.65 0.465 2.015 0.465 2.015 0.405 2.075 0.405 2.075 0.465 2.425 0.465 2.425 0.275 2.485 0.275 2.485 0.335 2.745 0.335 2.745 0.305 2.925 0.305 2.925 0.285 3.385 0.285 3.385 0.305 3.455 0.305 3.455 0.365 3.335 0.365 3.335 0.345 2.985 0.345 2.985 0.365 2.805 0.365 2.805 0.525 1.65 0.525 1.65 0.825 1.21 0.825 1.21 0.775 0.89 0.775 0.89 1.085 1.605 1.085 1.605 1.33 2.325 1.33 2.325 1.435 2.735 1.435 2.735 1.38 3.625 1.38 3.625 1.315 4.785 1.315 4.785 0.525 3.96 0.525 3.96 0.505 3.89 0.505 3.89 0.445 4.01 0.445 4.01 0.465 4.33 0.465 4.33 0.445 4.45 0.445 4.45 0.465 4.785 0.465 4.785 0.415 4.845 0.415 ;
      RECT 3.645 0.665 4.375 0.745 ;
      POLYGON 2.805 0.895 2.04 0.895 2.04 0.985 1.05 0.985 1.05 0.935 0.99 0.935 0.99 0.875 1.11 0.875 1.11 0.925 1.92 0.925 1.92 0.835 2.805 0.835 ;
      RECT 1.75 0.625 2.375 0.705 ;
      POLYGON 1.49 0.665 1.37 0.665 1.37 0.555 1.225 0.555 1.225 0.345 0.57 0.345 0.57 0.585 0.16 0.585 0.16 1.285 0.24 1.285 0.24 1.405 0.18 1.405 0.18 1.345 0.1 1.345 0.1 0.525 0.145 0.525 0.145 0.445 0.205 0.445 0.205 0.525 0.51 0.525 0.51 0.285 1.285 0.285 1.285 0.495 1.43 0.495 1.43 0.605 1.49 0.605 ;
      POLYGON 0.73 1.345 0.65 1.345 0.65 1.405 0.59 1.405 0.59 1.285 0.67 1.285 0.67 0.445 0.73 0.445 ;
  END
END OAI2BB2X4

MACRO OAI2BB2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI2BB2XL 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0395 LAYER Metal1 ;
    ANTENNADIFFAREA 1.03195 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 32.08333325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 258.8425925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.9 1.21 1.765 1.21 1.765 1.275 1.555 1.275 1.555 1.215 1.635 1.215 1.635 1.15 1.84 1.15 1.84 0.355 1.9 0.355 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.14 0.73 2.08 0.73 2.08 1.04 2 1.04 2 0.65 2.06 0.65 2.06 0.6 2.14 0.6 ;
    END
  END B0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.55 1.74 1.05 ;
    END
  END B1
  PIN A0N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.59 0.54 1.09 ;
    END
  END A0N
  PIN A1N
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.5 0.34 1 ;
    END
  END A1N
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.335 1.65 0.335 1.175 0.395 1.175 0.395 1.65 1.275 1.65 1.275 1.28 1.335 1.28 1.335 1.65 1.865 1.65 1.865 1.31 1.985 1.31 1.985 1.37 1.925 1.37 1.925 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 1.24 0.06 1.24 0.45 1.18 0.45 1.18 0.06 0.355 0.06 0.355 0.2 0.295 0.2 0.295 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.105 0.45 2.045 0.45 2.045 0.255 1.74 0.255 1.74 0.39 1.645 0.39 1.645 0.45 1.56 0.45 1.56 0.77 0.86 0.77 0.86 0.355 0.92 0.355 0.92 0.71 1.5 0.71 1.5 0.39 1.585 0.39 1.585 0.33 1.68 0.33 1.68 0.195 2.105 0.195 ;
      POLYGON 1.545 0.23 1.4 0.23 1.4 0.61 1.02 0.61 1.02 0.255 0.515 0.255 0.515 0.4 0.16 0.4 0.16 1.08 0.19 1.08 0.19 1.2 0.13 1.2 0.13 1.14 0.1 1.14 0.1 0.34 0.455 0.34 0.455 0.195 1.08 0.195 1.08 0.55 1.34 0.55 1.34 0.17 1.545 0.17 ;
      POLYGON 1.13 0.93 0.7 0.93 0.7 1.2 0.64 1.2 0.64 0.49 0.615 0.49 0.615 0.37 0.675 0.37 0.675 0.43 0.7 0.43 0.7 0.87 1.13 0.87 ;
  END
END OAI2BB2XL

MACRO OAI31X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.556825 LAYER Metal1 ;
    ANTENNADIFFAREA 0.7378 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.07 1.16 0.79 1.16 0.79 1.48 0.73 1.48 0.73 1.1 1.01 1.1 1.01 0.54 0.99 0.54 0.99 0.23 1.07 0.23 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.25 0.87 0.14 0.87 0.14 0.92 0.06 0.92 0.06 0.79 0.17 0.79 0.17 0.6 0.25 0.6 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.12820525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.6 0.94 1.02 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.6 0.74 1.04 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.245 1.65 0.245 1.09 0.305 1.09 0.305 1.65 0.935 1.65 0.935 1.24 0.995 1.24 0.995 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.65 0.06 0.65 0.32 0.53 0.32 0.53 0.06 0.205 0.06 0.205 0.47 0.145 0.47 0.145 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.83 0.5 0.35 0.5 0.35 0.23 0.41 0.23 0.41 0.435 0.765 0.435 0.765 0.23 0.83 0.23 ;
  END
END OAI31X1

MACRO OAI31X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X2 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.913925 LAYER Metal1 ;
    ANTENNADIFFAREA 1.5813 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.875 0.605 1.76 0.605 1.76 1.11 1.715 1.11 1.715 1.435 1.655 1.435 1.655 1.245 0.97 1.245 0.97 1.305 0.91 1.305 0.91 1.185 1.46 1.185 1.46 0.98 1.54 0.98 1.54 1.05 1.7 1.05 1.7 0.545 1.875 0.545 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.3 0.995 1.165 0.995 1.165 1.085 0.89 1.085 0.89 1.005 0.945 1.005 0.945 0.915 1.3 0.915 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.64102575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.235 0.815 0.74 0.815 0.74 0.92 0.66 0.92 0.66 0.815 0.495 0.815 0.495 0.755 1.235 0.755 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.051282 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 0.82 1.4 0.82 1.4 0.655 0.395 0.655 0.395 0.795 0.335 0.795 0.335 0.595 1.46 0.595 1.46 0.6 1.54 0.6 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.705 1.94 1.205 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.29 1.65 0.29 1.045 0.35 1.045 0.35 1.65 1.42 1.65 1.42 1.345 1.54 1.345 1.54 1.405 1.48 1.405 1.48 1.65 1.86 1.65 1.86 1.305 1.92 1.305 1.92 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 1.335 0.06 1.335 0.16 1.395 0.16 1.395 0.22 1.275 0.22 1.275 0.06 0.865 0.06 0.865 0.16 0.925 0.16 0.925 0.22 0.805 0.22 0.805 0.06 0.395 0.06 0.395 0.16 0.455 0.16 0.455 0.22 0.335 0.22 0.335 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.05 0.495 1.99 0.495 1.99 0.435 1.6 0.435 1.6 0.495 0.1 0.495 0.1 0.435 1.54 0.435 1.54 0.375 2.05 0.375 ;
  END
END OAI31X2

MACRO OAI31X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31X4 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.720375 LAYER Metal1 ;
    ANTENNADIFFAREA 3.0637 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.675 0.545 3.6 0.545 3.6 0.595 3.12 0.595 3.12 0.98 3.14 0.98 3.14 1.05 3.485 1.05 3.485 1.015 3.545 1.015 3.545 1.405 3.485 1.405 3.485 1.11 3.135 1.11 3.135 1.405 3.075 1.405 3.075 1.185 2.225 1.185 2.225 1.405 2.165 1.405 2.165 1.185 0.975 1.185 0.975 1.405 0.915 1.405 0.915 1.125 3.06 1.125 3.06 0.485 3.265 0.485 3.265 0.535 3.54 0.535 3.54 0.485 3.675 0.485 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.705 0.895 3.425 0.895 3.425 0.88 3.22 0.88 3.22 0.8 3.705 0.8 ;
    END
  END B0
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.65384625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.82 1.025 0.605 1.025 0.605 0.935 0.235 0.935 0.235 0.815 0.365 0.815 0.365 0.875 0.665 0.875 0.665 0.965 1.425 0.965 1.425 0.885 1.545 0.885 1.545 0.965 2.76 0.965 2.76 0.855 2.82 0.855 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.9102565 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.565 0.745 2.32 0.745 2.32 0.865 1.645 0.865 1.645 0.785 1.325 0.785 1.325 0.865 0.765 0.865 0.765 0.715 0.445 0.715 0.445 0.655 0.825 0.655 0.825 0.805 1.265 0.805 1.265 0.725 1.705 0.725 1.705 0.805 2.26 0.805 2.26 0.6 2.34 0.6 2.34 0.625 2.565 0.625 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.6153845 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.115 0.705 1.805 0.705 1.805 0.625 1.165 0.625 1.165 0.705 0.925 0.705 0.925 0.645 1.035 0.645 1.035 0.625 1.105 0.625 1.105 0.565 1.865 0.565 1.865 0.645 2.115 0.645 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 0 1.77 0 1.65 0.24 1.65 0.24 1.035 0.3 1.035 0.3 1.65 1.49 1.65 1.49 1.285 1.55 1.285 1.55 1.65 2.825 1.65 2.825 1.285 2.885 1.285 2.885 1.65 3.28 1.65 3.28 1.285 3.34 1.285 3.34 1.65 3.69 1.65 3.69 1.015 3.75 1.015 3.75 1.65 4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 2.695 0.06 2.695 0.16 2.755 0.16 2.755 0.22 2.635 0.22 2.635 0.06 2.225 0.06 2.225 0.16 2.285 0.16 2.285 0.22 2.165 0.22 2.165 0.06 1.755 0.06 1.755 0.16 1.815 0.16 1.815 0.22 1.695 0.22 1.695 0.06 1.285 0.06 1.285 0.16 1.345 0.16 1.345 0.22 1.225 0.22 1.225 0.06 0.815 0.06 0.815 0.16 0.875 0.16 0.875 0.22 0.755 0.22 0.755 0.06 0.345 0.06 0.345 0.16 0.405 0.16 0.405 0.22 0.285 0.22 0.285 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.85 0.435 3.79 0.435 3.79 0.375 3.44 0.375 3.44 0.435 3.38 0.435 3.38 0.375 2.96 0.375 2.96 0.435 0.05 0.435 0.05 0.375 2.9 0.375 2.9 0.315 3.85 0.315 ;
  END
END OAI31X4

MACRO OAI31XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI31XL 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5751 LAYER Metal1 ;
    ANTENNADIFFAREA 0.6264 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 1.11 0.9 1.11 0.9 1.27 0.855 1.27 0.855 1.33 0.795 1.33 0.795 1.21 0.84 1.21 0.84 0.98 1.08 0.98 1.08 0.255 1.14 0.255 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END A1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.6 0.14 1.1 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.98 0.88 0.86 0.88 0.86 0.6 0.9 0.6 0.9 0.42 0.98 0.42 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.61 0.74 1.11 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.23 1.65 0.23 1.21 0.29 1.21 0.29 1.65 1 1.65 1 1.21 1.06 1.21 1.06 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 0.6 0.06 0.6 0.35 0.54 0.35 0.54 0.06 0.13 0.06 0.13 0.35 0.07 0.35 0.07 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.835 0.32 0.76 0.32 0.76 0.51 0.335 0.51 0.335 0.255 0.395 0.255 0.395 0.45 0.7 0.45 0.7 0.26 0.835 0.26 ;
  END
END OAI31XL

MACRO OAI32X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.56815 LAYER Metal1 ;
    ANTENNADIFFAREA 0.92035 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.95 0.73 0.745 0.73 0.745 1.48 0.665 1.48 0.665 0.67 0.89 0.67 0.89 0.32 0.95 0.32 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.79487175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.3 0.695 0.14 0.695 0.14 0.94 0.06 0.94 0.06 0.615 0.3 0.615 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20512825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.365 0.945 0.34 0.945 0.34 1.3 0.26 1.3 0.26 0.8 0.365 0.8 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.815 0.81 0.96 0.955 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.79487175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.585 0.83 0.54 0.83 0.54 1.13 0.46 1.13 0.46 0.745 0.505 0.745 0.505 0.69 0.585 0.69 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.71794875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.17 0.705 1.14 0.705 1.14 0.925 1.05 0.925 1.05 0.705 1.02 0.705 1.02 0.615 1.17 0.615 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1 0.13 1 0.13 1.65 1.06 1.65 1.06 1 1.12 1 1.12 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 0.51 0.06 0.51 0.33 0.57 0.33 0.57 0.39 0.45 0.39 0.45 0.06 0.13 0.06 0.13 0.54 0.07 0.54 0.07 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.155 0.54 1.095 0.54 1.095 0.25 0.745 0.25 0.745 0.55 0.275 0.55 0.275 0.3 0.335 0.3 0.335 0.49 0.685 0.49 0.685 0.185 1.155 0.185 ;
  END
END OAI32X1

MACRO OAI32X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X2 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1063 LAYER Metal1 ;
    ANTENNADIFFAREA 1.85355 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.26 0.515 2.185 0.515 2.185 0.565 1.5 0.565 1.5 1.245 1.925 1.245 1.925 1.365 1.865 1.365 1.865 1.305 1.44 1.305 1.44 1.085 0.87 1.085 0.87 1.365 0.81 1.365 0.81 1.025 1.235 1.025 1.235 1.005 1.44 1.005 1.44 0.505 1.73 0.505 1.73 0.455 1.85 0.455 1.85 0.505 2.125 0.505 2.125 0.455 2.26 0.455 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.76 0.925 0.54 0.925 0.54 1.125 0.46 1.125 0.46 0.845 0.76 0.845 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.84615375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.16 0.785 0.94 0.785 0.94 0.92 0.86 0.92 0.86 0.745 0.47 0.745 0.47 0.665 1.16 0.665 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.1 0.905 1.94 0.905 1.94 1.145 1.86 1.145 1.86 0.905 1.84 0.905 1.84 0.825 2.1 0.825 ;
    END
  END B1
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.73 1.26 0.73 1.26 0.565 0.295 0.565 0.295 0.73 0.235 0.73 0.235 0.505 1.34 0.505 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.897436 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.3 0.725 1.74 0.725 1.74 0.92 1.66 0.92 1.66 0.725 1.6 0.725 1.6 0.665 2.3 0.665 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 1.77 0 1.77 0 1.65 0.265 1.65 0.265 0.975 0.325 0.975 0.325 1.65 1.42 1.65 1.42 1.405 1.54 1.405 1.54 1.465 1.48 1.465 1.48 1.65 2.2 1.65 2.2 0.975 2.26 0.975 2.26 1.65 2.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 0.06 1.3 0.06 1.3 0.16 1.36 0.16 1.36 0.22 1.24 0.22 1.24 0.06 0.83 0.06 0.83 0.16 0.89 0.16 0.89 0.22 0.77 0.22 0.77 0.06 0.36 0.06 0.36 0.16 0.42 0.16 0.42 0.22 0.3 0.22 0.3 0.06 0 0.06 0 -0.06 2.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.435 0.405 2.375 0.405 2.375 0.345 2.025 0.345 2.025 0.405 1.965 0.405 1.965 0.345 1.565 0.345 1.565 0.405 0.065 0.405 0.065 0.345 1.505 0.345 1.505 0.285 2.435 0.285 ;
  END
END OAI32X2

MACRO OAI32X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32X4 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9854 LAYER Metal1 ;
    ANTENNADIFFAREA 3.51835 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.415 0.545 4.34 0.545 4.34 0.595 3.125 0.595 3.125 0.745 2.915 0.745 2.915 1.155 3.93 1.155 3.93 1.275 3.87 1.275 3.87 1.215 3.31 1.215 3.31 1.275 3.25 1.275 3.25 1.215 2.565 1.215 2.565 1.275 2.435 1.275 2.435 1.215 2.215 1.215 2.215 1.275 2.155 1.275 2.155 1.215 0.965 1.215 0.965 1.275 0.905 1.275 0.905 1.155 2.855 1.155 2.855 0.685 3.065 0.685 3.065 0.485 3.185 0.485 3.185 0.535 3.475 0.535 3.475 0.485 3.595 0.485 3.595 0.535 3.885 0.535 3.885 0.485 4.005 0.485 4.005 0.535 4.28 0.535 4.28 0.485 4.415 0.485 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.71794875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.755 1.055 0.32 1.055 0.32 0.895 0.235 0.895 0.235 0.815 0.38 0.815 0.38 0.995 1.425 0.995 1.425 0.885 1.545 0.885 1.545 0.995 2.695 0.995 2.695 0.855 2.755 0.855 ;
    END
  END A0
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.74358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.34 0.92 4.175 0.92 4.175 1.055 3.015 1.055 3.015 0.845 3.075 0.845 3.075 0.995 3.595 0.995 3.595 0.885 3.715 0.885 3.715 0.995 4.115 0.995 4.115 0.855 4.26 0.855 4.26 0.79 4.34 0.79 ;
    END
  END B0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.1153845 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.585 0.895 1.8 0.895 1.8 0.785 1.325 0.785 1.325 0.875 0.765 0.875 0.765 0.895 0.635 0.895 0.635 0.875 0.48 0.875 0.48 0.815 1.265 0.815 1.265 0.725 1.86 0.725 1.86 0.835 2.585 0.835 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.25641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.005 0.895 3.835 0.895 3.835 0.785 3.295 0.785 3.295 0.725 3.895 0.725 3.895 0.775 4.005 0.775 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.6153845 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.075 0.735 2.015 0.735 2.015 0.625 1.165 0.625 1.165 0.705 0.915 0.705 0.915 0.645 1.035 0.645 1.035 0.625 1.105 0.625 1.105 0.565 2.075 0.565 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.275 1.65 0.275 1.285 0.335 1.285 0.335 1.65 1.565 1.65 1.565 1.315 1.685 1.315 1.685 1.375 1.625 1.375 1.625 1.65 2.835 1.65 2.835 1.375 2.955 1.375 2.955 1.435 2.895 1.435 2.895 1.65 3.53 1.65 3.53 1.315 3.65 1.315 3.65 1.375 3.59 1.375 3.59 1.65 4.18 1.65 4.18 1.285 4.24 1.285 4.24 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 2.685 0.06 2.685 0.16 2.745 0.16 2.745 0.22 2.625 0.22 2.625 0.06 2.215 0.06 2.215 0.16 2.275 0.16 2.275 0.22 2.155 0.22 2.155 0.06 1.745 0.06 1.745 0.16 1.805 0.16 1.805 0.22 1.685 0.22 1.685 0.06 1.275 0.06 1.275 0.16 1.335 0.16 1.335 0.22 1.215 0.22 1.215 0.06 0.805 0.06 0.805 0.16 0.865 0.16 0.865 0.22 0.745 0.22 0.745 0.06 0.335 0.06 0.335 0.16 0.395 0.16 0.395 0.22 0.275 0.22 0.275 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.59 0.435 4.53 0.435 4.53 0.375 4.18 0.375 4.18 0.435 4.12 0.435 4.12 0.375 3.77 0.375 3.77 0.435 3.71 0.435 3.71 0.375 3.36 0.375 3.36 0.435 3.3 0.435 3.3 0.375 2.95 0.375 2.95 0.435 0.04 0.435 0.04 0.375 2.89 0.375 2.89 0.315 4.59 0.315 ;
  END
END OAI32X4

MACRO OAI32XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI32XL 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6456 LAYER Metal1 ;
    ANTENNADIFFAREA 0.841625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.3 0.8 1.165 0.8 1.165 1.235 1.105 1.235 1.105 1.085 1.035 1.085 1.035 1.005 1.105 1.005 1.105 0.74 1.24 0.74 1.24 0.415 1.3 0.415 ;
    END
  END Y
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.61 0.34 1.11 ;
    END
  END A0
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 1.27 0.48 1.27 0.48 0.92 0.46 0.92 0.46 0.79 0.56 0.79 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 1.11 1.265 1.11 1.265 0.9 1.345 0.9 1.345 1.03 1.46 1.03 1.46 0.935 1.54 0.935 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.005 0.82 0.74 0.82 0.74 0.975 0.66 0.975 0.66 0.74 1.005 0.74 ;
    END
  END A2
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 0.92 1.66 0.92 1.66 0.8 1.425 0.8 1.425 0.655 1.505 0.655 1.505 0.72 1.74 0.72 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.235 1.65 0.235 1.21 0.295 1.21 0.295 1.65 1.5 1.65 1.5 1.21 1.56 1.21 1.56 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 0.675 0.06 0.675 0.42 0.735 0.42 0.735 0.48 0.615 0.48 0.615 0.06 0.295 0.06 0.295 0.51 0.235 0.51 0.235 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.505 0.51 1.445 0.51 1.445 0.315 0.91 0.315 0.91 0.64 0.44 0.64 0.44 0.415 0.5 0.415 0.5 0.58 0.85 0.58 0.85 0.255 1.505 0.255 ;
  END
END OAI32XL

MACRO OAI33X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X1 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7087 LAYER Metal1 ;
    ANTENNADIFFAREA 1.02555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 1.27 0.845 1.27 0.845 1.46 0.785 1.46 0.785 1.21 1.44 1.21 1.44 0.51 0.99 0.51 0.99 0.37 1.05 0.37 1.05 0.45 1.4 0.45 1.4 0.37 1.5 0.37 1.5 0.98 1.54 0.98 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.86 0.61 0.94 1.11 ;
    END
  END B2
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.61 0.34 1.11 ;
    END
  END A0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.61 0.74 1.11 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.61 1.14 1.11 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.61 1.34 1.11 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.24 1.65 0.24 1.21 0.3 1.21 0.3 1.65 1.265 1.65 1.265 1.37 1.385 1.37 1.385 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 0.61 0.06 0.61 0.35 0.55 0.35 0.55 0.06 0.2 0.06 0.2 0.35 0.14 0.35 0.14 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.255 0.35 1.195 0.35 1.195 0.27 0.815 0.27 0.815 0.51 0.345 0.51 0.345 0.37 0.405 0.37 0.405 0.45 0.755 0.45 0.755 0.21 1.255 0.21 ;
  END
END OAI33X1

MACRO OAI33X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X2 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.05895 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.76844775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.03 1.065 3.165 1.065 3.165 1.085 3.03 1.085 3.03 1.065 2.84 1.065 2.84 1.005 3.97 1.005 3.97 0.945 4.03 0.945 ;
    END
  END B0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.05895 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.01526725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.235 1.085 2.035 1.085 2.035 1.055 0.75 1.055 0.75 0.995 2.235 0.995 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.05895 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.50636125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.87 0.905 2.74 0.905 2.74 1.11 2.66 1.11 2.66 0.98 2.68 0.98 2.68 0.845 3.87 0.845 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.05895 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.7862595 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.935 0.895 1.635 0.895 1.635 0.875 0.485 0.875 0.485 0.815 1.935 0.815 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.05895 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.557252 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.71 0.745 2.54 0.745 2.54 0.92 2.46 0.92 2.46 0.685 3.71 0.685 ;
    END
  END B2
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.05895 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.3867685 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.5 0.705 0.325 0.705 0.325 0.645 0.435 0.645 0.435 0.625 0.565 0.625 0.565 0.645 1.5 0.645 ;
    END
  END A0
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.96115 LAYER Metal1 ;
    ANTENNADIFFAREA 2.502175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.295 0.505 4.25 0.505 4.25 0.635 4.19 0.635 4.19 1.27 0.835 1.27 0.835 1.21 4.13 1.21 4.13 0.635 3.81 0.635 3.81 0.585 2.535 0.585 2.535 0.515 2.435 0.515 2.435 0.435 2.475 0.435 2.475 0.415 2.595 0.415 2.595 0.525 2.915 0.525 2.915 0.415 3.035 0.415 3.035 0.525 3.355 0.525 3.355 0.415 3.475 0.415 3.475 0.525 3.795 0.525 3.795 0.415 3.915 0.415 3.915 0.475 3.87 0.475 3.87 0.575 4.19 0.575 4.19 0.445 4.235 0.445 4.235 0.385 4.295 0.385 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.28 1.65 0.28 1.28 0.34 1.28 0.34 1.65 1.335 1.65 1.335 1.37 1.455 1.37 1.455 1.43 1.395 1.43 1.395 1.65 2.935 1.65 2.935 1.37 3.055 1.37 3.055 1.43 2.995 1.43 2.995 1.65 4.045 1.65 4.045 1.37 4.165 1.37 4.165 1.43 4.105 1.43 4.105 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 2.07 0.06 2.07 0.305 2.13 0.305 2.13 0.365 2.01 0.365 2.01 0.06 1.6 0.06 1.6 0.305 1.66 0.305 1.66 0.365 1.54 0.365 1.54 0.06 1.13 0.06 1.13 0.305 1.19 0.305 1.19 0.365 1.07 0.365 1.07 0.06 0.65 0.06 0.65 0.305 0.71 0.305 0.71 0.365 0.59 0.365 0.59 0.06 0.24 0.06 0.24 0.445 0.18 0.445 0.18 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.09 0.455 4.03 0.455 4.03 0.315 3.695 0.315 3.695 0.425 3.575 0.425 3.575 0.315 3.255 0.315 3.255 0.42 3.135 0.42 3.135 0.315 2.815 0.315 2.815 0.42 2.695 0.42 2.695 0.315 2.335 0.315 2.335 0.525 0.385 0.525 0.385 0.38 0.445 0.38 0.445 0.465 0.855 0.465 0.855 0.38 0.915 0.38 0.915 0.465 1.335 0.465 1.335 0.38 1.395 0.38 1.395 0.465 1.805 0.465 1.805 0.38 1.865 0.38 1.865 0.465 2.275 0.465 2.275 0.255 4.09 0.255 ;
  END
END OAI33X2

MACRO OAI33X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33X4 0 0 ;
  SIZE 5.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.924 LAYER Metal1 ;
    ANTENNADIFFAREA 4.0726 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.21 0.535 5.135 0.535 5.135 0.585 3.09 0.585 3.09 0.715 2.165 0.715 2.165 0.995 3.745 0.995 3.745 1.185 3.685 1.185 3.685 1.055 3.325 1.055 3.325 1.185 3.265 1.185 3.265 1.055 2.915 1.055 2.915 1.345 2.855 1.345 2.855 1.055 2.495 1.055 2.495 1.185 2.435 1.185 2.435 1.055 2.085 1.055 2.085 1.185 2.025 1.185 2.025 0.995 2.105 0.995 2.105 0.895 2.035 0.895 2.035 0.815 2.105 0.815 2.105 0.655 3.03 0.655 3.03 0.475 3.15 0.475 3.15 0.525 3.45 0.525 3.45 0.475 3.57 0.475 3.57 0.525 3.86 0.525 3.86 0.475 3.98 0.475 3.98 0.525 4.27 0.525 4.27 0.475 4.39 0.475 4.39 0.525 4.68 0.525 4.68 0.475 4.8 0.475 4.8 0.525 5.075 0.525 5.075 0.475 5.21 0.475 ;
    END
  END Y
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.79487175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.34 0.895 4.85 0.895 4.85 0.685 4.93 0.685 4.93 0.815 5.34 0.815 ;
    END
  END B0
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.14 0.815 3.64 0.895 ;
    END
  END B2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.9358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 0.92 1.66 0.92 1.66 0.895 1.25 0.895 1.25 0.815 1.66 0.815 1.66 0.655 1.74 0.655 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.4871795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.265 0.815 2.765 0.895 ;
    END
  END A2
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.82051275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 0.92 0.495 0.92 0.495 0.84 0.86 0.84 0.86 0.655 0.94 0.655 ;
    END
  END A0
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.67948725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.455 0.895 4.01 0.895 4.01 0.685 4.165 0.685 4.165 0.815 4.455 0.815 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 1.77 0 1.77 0 1.65 0.385 1.65 0.385 1.265 0.445 1.265 0.445 1.65 0.795 1.65 0.795 1.265 0.855 1.265 0.855 1.65 4.915 1.65 4.915 1.255 4.975 1.255 4.975 1.65 5.325 1.65 5.325 1.255 5.385 1.255 5.385 1.65 5.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 0.06 2.68 0.06 2.68 0.335 2.74 0.335 2.74 0.395 2.62 0.395 2.62 0.06 2.26 0.06 2.26 0.335 2.32 0.335 2.32 0.395 2.2 0.395 2.2 0.06 1.85 0.06 1.85 0.335 1.91 0.335 1.91 0.395 1.79 0.395 1.79 0.06 1.44 0.06 1.44 0.335 1.5 0.335 1.5 0.395 1.38 0.395 1.38 0.06 1.03 0.06 1.03 0.335 1.09 0.335 1.09 0.395 0.97 0.395 0.97 0.06 0.62 0.06 0.62 0.335 0.68 0.335 0.68 0.395 0.56 0.395 0.56 0.06 0 0.06 0 -0.06 5.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.59 1.375 5.53 1.375 5.53 1.055 5.18 1.055 5.18 1.375 5.12 1.375 5.12 1.055 4.77 1.055 4.77 1.375 4.71 1.375 4.71 1.055 4.36 1.055 4.36 1.115 4.3 1.115 4.3 1.055 3.95 1.055 3.95 1.115 3.89 1.115 3.89 0.995 5.59 0.995 ;
      POLYGON 5.385 0.425 5.325 0.425 5.325 0.365 4.975 0.365 4.975 0.425 4.915 0.425 4.915 0.365 4.565 0.365 4.565 0.425 4.505 0.425 4.505 0.365 4.155 0.365 4.155 0.425 4.095 0.425 4.095 0.365 3.745 0.365 3.745 0.425 3.685 0.425 3.685 0.365 3.325 0.365 3.325 0.425 3.265 0.425 3.265 0.365 2.915 0.365 2.915 0.555 0.385 0.555 0.385 0.435 0.445 0.435 0.445 0.495 0.795 0.495 0.795 0.435 0.855 0.435 0.855 0.495 1.205 0.495 1.205 0.435 1.265 0.435 1.265 0.495 1.615 0.495 1.615 0.435 1.675 0.435 1.675 0.495 2.025 0.495 2.025 0.435 2.085 0.435 2.085 0.495 2.435 0.495 2.435 0.435 2.495 0.435 2.495 0.495 2.855 0.495 2.855 0.305 5.385 0.305 ;
      POLYGON 4.565 1.345 3.06 1.345 3.06 1.225 3.12 1.225 3.12 1.285 3.48 1.285 3.48 1.225 3.54 1.225 3.54 1.285 4.095 1.285 4.095 1.225 4.155 1.225 4.155 1.285 4.505 1.285 4.505 1.225 4.565 1.225 ;
      POLYGON 2.71 1.345 1.205 1.345 1.205 1.225 1.265 1.225 1.265 1.285 1.615 1.285 1.615 1.225 1.675 1.225 1.675 1.285 2.23 1.285 2.23 1.225 2.29 1.225 2.29 1.285 2.65 1.285 2.65 1.225 2.71 1.225 ;
      POLYGON 1.88 1.14 1.82 1.14 1.82 1.08 1.47 1.08 1.47 1.14 1.41 1.14 1.41 1.08 1.06 1.08 1.06 1.385 1 1.385 1 1.08 0.65 1.08 0.65 1.385 0.59 1.385 0.59 1.08 0.24 1.08 0.24 1.385 0.18 1.385 0.18 1.02 1.88 1.02 ;
  END
END OAI33X4

MACRO OAI33XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI33XL 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.775625 LAYER Metal1 ;
    ANTENNADIFFAREA 0.8613 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 1.245 1.025 1.245 1.025 1.37 0.965 1.37 0.965 1.185 1.66 1.185 1.66 0.98 1.68 0.98 1.68 0.485 1.2 0.485 1.2 0.35 1.14 0.35 1.14 0.29 1.26 0.29 1.26 0.425 1.595 0.425 1.595 0.26 1.74 0.26 ;
    END
  END Y
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.745 0.54 1.245 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.13 1.085 0.86 1.085 0.86 0.775 0.94 0.775 0.94 1.005 1.13 1.005 ;
    END
  END B2
  PIN A0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.32 0.92 0.22 0.92 0.22 0.73 0.06 0.73 0.06 0.6 0.14 0.6 0.14 0.65 0.32 0.65 ;
    END
  END A0
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.79 0.74 1.29 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.585 1.34 1.085 ;
    END
  END B1
  PIN B0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 1.065 1.46 1.065 1.46 0.705 1.44 0.705 1.44 0.585 1.52 0.585 1.52 0.6 1.54 0.6 ;
    END
  END B0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.245 1.65 0.245 1.345 0.305 1.345 0.305 1.65 1.515 1.65 1.515 1.345 1.575 1.345 1.575 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 0.615 0.06 0.615 0.355 0.555 0.355 0.555 0.06 0.205 0.06 0.205 0.355 0.145 0.355 0.145 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.48 0.325 1.36 0.325 1.36 0.22 0.85 0.22 0.85 0.515 0.35 0.515 0.35 0.26 0.41 0.26 0.41 0.455 0.79 0.455 0.79 0.16 1.42 0.16 1.42 0.265 1.48 0.265 ;
  END
END OAI33XL

MACRO OR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X1 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3636 LAYER Metal1 ;
    ANTENNADIFFAREA 0.50205 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.43076925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 102.6153845 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.75 0.94 0.73 0.94 0.73 1.29 0.67 1.29 0.67 0.895 0.66 0.895 0.66 0.815 0.67 0.815 0.67 0.375 0.73 0.375 0.73 0.595 0.75 0.595 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.27777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.45 0.82 0.39 0.82 0.39 1.055 0.34 1.055 0.34 1.125 0.26 1.125 0.26 0.98 0.32 0.98 0.32 0.76 0.45 0.76 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.04 0.58 0.14 0.8 ;
    END
  END B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 0.06 0.495 0.06 0.495 0.51 0.555 0.51 0.555 0.58 0.435 0.58 0.435 0.06 0.185 0.06 0.185 0.3 0.065 0.3 0.065 0.06 0 0.06 0 -0.06 0.8 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.77 0 1.77 0 1.65 0.465 1.65 0.465 0.91 0.525 0.91 0.525 1.65 0.8 1.65 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 0.595 0.81 0.535 0.81 0.535 0.7 0.26 0.7 0.26 0.92 0.185 0.92 0.185 1.025 0.125 1.025 0.125 0.86 0.2 0.86 0.2 0.63 0.26 0.63 0.26 0.505 0.32 0.505 0.32 0.64 0.595 0.64 ;
  END
END OR2X1

MACRO OR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X2 0 0 ;
  SIZE 1 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.442175 LAYER Metal1 ;
    ANTENNADIFFAREA 0.674775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.558547 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 58.025641 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 0.925 0.735 0.925 0.735 1.34 0.675 1.34 0.675 0.925 0.66 0.925 0.66 0.59 0.675 0.59 0.675 0.385 0.735 0.385 0.735 0.59 0.74 0.59 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.83333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.445 0.85 0.395 0.85 0.395 0.99 0.34 0.99 0.34 1.13 0.26 1.13 0.26 0.91 0.32 0.91 0.32 0.73 0.445 0.73 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.045 0.41 0.14 0.72 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.77 0 1.77 0 1.65 0.47 1.65 0.47 0.98 0.53 0.98 0.53 1.65 0.81 1.65 0.81 1.51 0.93 1.51 0.93 1.65 1 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.06 0.93 0.06 0.93 0.215 0.805 0.215 0.805 0.06 0.5 0.06 0.5 0.445 0.56 0.445 0.56 0.505 0.44 0.505 0.44 0.06 0.17 0.06 0.17 0.245 0.04 0.245 0.04 0.06 0 0.06 0 -0.06 1 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.59 0.815 0.53 0.815 0.53 0.665 0.26 0.665 0.26 0.845 0.19 0.845 0.19 1.075 0.13 1.075 0.13 0.78 0.2 0.78 0.2 0.605 0.235 0.605 0.235 0.44 0.295 0.44 0.295 0.605 0.59 0.605 ;
  END
END OR2X2

MACRO OR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X4 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.93175 LAYER Metal1 ;
    ANTENNADIFFAREA 1.0665 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.96367525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 62.25641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 0.73 1.305 0.73 1.305 1.075 1.245 1.075 1.245 1.405 1.185 1.405 1.185 1.015 1.245 1.015 1.245 0.915 0.82 0.915 0.82 1.405 0.76 1.405 0.76 0.855 1.245 0.855 1.245 0.73 1.235 0.73 1.235 0.59 0.76 0.59 0.76 0.23 0.82 0.23 0.82 0.53 1.185 0.53 1.185 0.23 1.245 0.23 1.245 0.53 1.305 0.53 1.305 0.6 1.365 0.6 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.12820525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.565 1.085 0.435 1.085 0.435 1.005 0.445 1.005 0.445 0.715 0.54 0.715 0.54 1.005 0.565 1.005 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.12820525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.22 0.925 0.06 0.925 0.06 0.785 0.14 0.785 0.14 0.585 0.22 0.585 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.54 1.65 0.54 1.165 0.6 1.165 0.6 1.65 0.965 1.65 0.965 1.015 1.025 1.015 1.025 1.65 1.39 1.65 1.39 1.015 1.45 1.015 1.45 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.45 0.06 1.45 0.47 1.39 0.47 1.39 0.06 1.04 0.06 1.04 0.47 0.98 0.47 0.98 0.06 0.6 0.06 0.6 0.49 0.54 0.49 0.54 0.06 0.19 0.06 0.19 0.49 0.13 0.49 0.13 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.145 0.715 0.635 0.715 0.635 0.655 0.355 0.655 0.355 1.405 0.23 1.405 0.23 1.015 0.29 1.015 0.29 0.585 0.335 0.585 0.335 0.23 0.395 0.23 0.395 0.585 0.7 0.585 0.7 0.655 1.145 0.655 ;
  END
END OR2X4

MACRO OR2X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X6 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2883 LAYER Metal1 ;
    ANTENNADIFFAREA 1.6252 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.34074075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 58.4957265 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.165 0.73 1.945 0.73 1.945 0.96 2.005 0.96 2.005 1.43 1.945 1.43 1.945 1.02 1.595 1.02 1.595 1.43 1.535 1.43 1.535 1.02 1.185 1.02 1.185 1.43 1.125 1.43 1.125 0.96 1.86 0.96 1.86 0.72 1.125 0.72 1.125 0.35 1.185 0.35 1.185 0.66 1.535 0.66 1.535 0.35 1.595 0.35 1.595 0.66 1.945 0.66 1.945 0.35 2.005 0.35 2.005 0.6 2.165 0.6 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.71794875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.43 0.91 0.565 1.11 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.87179475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.865 0.84 0.26 0.84 0.26 0.925 0.06 0.925 0.06 0.78 0.865 0.78 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.2 1.65 0.2 1.04 0.26 1.04 0.26 1.65 0.85 1.65 0.85 1.07 0.91 1.07 0.91 1.65 1.33 1.65 1.33 1.12 1.39 1.12 1.39 1.65 1.74 1.65 1.74 1.12 1.8 1.12 1.8 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 1.8 0.06 1.8 0.59 1.74 0.59 1.74 0.06 1.39 0.06 1.39 0.59 1.33 0.59 1.33 0.06 0.965 0.06 0.965 0.59 0.905 0.59 0.905 0.06 0.555 0.06 0.555 0.59 0.495 0.59 0.495 0.06 0.13 0.06 0.13 0.59 0.07 0.59 0.07 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.69 0.84 1.025 0.84 1.025 0.97 0.725 0.97 0.725 1.245 0.6 1.245 0.6 1.43 0.54 1.43 0.54 1.185 0.665 1.185 0.665 0.91 0.965 0.91 0.965 0.72 0.29 0.72 0.29 0.35 0.35 0.35 0.35 0.66 0.7 0.66 0.7 0.35 0.76 0.35 0.76 0.66 1.025 0.66 1.025 0.78 1.69 0.78 ;
  END
END OR2X6

MACRO OR2X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2X8 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 0.06 2.21 0.06 2.21 0.59 2.15 0.59 2.15 0.06 1.8 0.06 1.8 0.59 1.74 0.59 1.74 0.06 1.39 0.06 1.39 0.59 1.33 0.59 1.33 0.06 0.965 0.06 0.965 0.59 0.905 0.59 0.905 0.06 0.555 0.06 0.555 0.59 0.495 0.59 0.495 0.06 0.13 0.06 0.13 0.59 0.07 0.59 0.07 0.06 0 0.06 0 -0.06 2.6 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 1.77 0 1.77 0 1.65 0.2 1.65 0.2 1.04 0.26 1.04 0.26 1.65 0.85 1.65 0.85 1.07 0.91 1.07 0.91 1.65 1.33 1.65 1.33 1.12 1.39 1.12 1.39 1.65 1.74 1.65 1.74 1.12 1.8 1.12 1.8 1.65 2.15 1.65 2.15 1.12 2.21 1.12 2.21 1.65 2.6 1.65 ;
    END
  END VDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.84615375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.865 0.84 0.26 0.84 0.26 0.92 0.06 0.92 0.06 0.78 0.865 0.78 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 1.74358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.43 0.91 0.565 1.115 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.56275 LAYER Metal1 ;
    ANTENNADIFFAREA 1.9348 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.23625 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.61481475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 53.015873 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.54 0.73 2.355 0.73 2.355 0.96 2.415 0.96 2.415 1.43 2.355 1.43 2.355 1.02 2.005 1.02 2.005 1.43 1.945 1.43 1.945 1.02 1.595 1.02 1.595 1.43 1.535 1.43 1.535 1.02 1.185 1.02 1.185 1.43 1.125 1.43 1.125 0.96 2.26 0.96 2.26 0.72 1.125 0.72 1.125 0.35 1.185 0.35 1.185 0.66 1.535 0.66 1.535 0.35 1.595 0.35 1.595 0.66 1.945 0.66 1.945 0.35 2.005 0.35 2.005 0.66 2.355 0.66 2.355 0.35 2.415 0.35 2.415 0.6 2.54 0.6 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      POLYGON 2.1 0.84 1.025 0.84 1.025 0.97 0.725 0.97 0.725 1.25 0.6 1.25 0.6 1.43 0.54 1.43 0.54 1.19 0.665 1.19 0.665 0.91 0.965 0.91 0.965 0.72 0.29 0.72 0.29 0.35 0.35 0.35 0.35 0.66 0.7 0.66 0.7 0.35 0.76 0.35 0.76 0.66 1.025 0.66 1.025 0.78 2.1 0.78 ;
  END
END OR2X8

MACRO OR2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2XL 0 0 ;
  SIZE 0.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3447 LAYER Metal1 ;
    ANTENNADIFFAREA 0.44405 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 21.27777775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 163.14814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.725 1.085 0.645 1.085 0.645 0.79 0.655 0.79 0.655 0.435 0.725 0.435 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.12962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.545 0.995 0.465 0.995 0.465 0.91 0.365 0.91 0.365 0.79 0.545 0.79 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.388889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.055 0.63 0.135 0.895 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.77 0 1.77 0 1.65 0.44 1.65 0.44 1.06 0.5 1.06 0.5 1.65 0.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 0.06 0.56 0.06 0.56 0.24 0.44 0.24 0.44 0.06 0.175 0.06 0.175 0.24 0.04 0.24 0.04 0.06 0 0.06 0 -0.06 0.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.575 0.73 0.515 0.73 0.515 0.665 0.295 0.665 0.295 1.12 0.1 1.12 0.1 1.06 0.235 1.06 0.235 0.41 0.295 0.41 0.295 0.605 0.575 0.605 ;
  END
END OR2XL

MACRO OR3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.50955 LAYER Metal1 ;
    ANTENNADIFFAREA 0.6544 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 17.42051275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 143.076923 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.14 0.555 1.015 0.555 1.015 1.3 0.935 1.3 0.935 0.325 1.015 0.325 1.015 0.41 1.14 0.41 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.68518525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 0.92 0.605 0.92 0.605 0.64 0.685 0.64 0.685 0.785 0.74 0.785 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.22222225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.835 0.375 1.11 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.27777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.035 0.625 0.18 0.765 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.73 1.65 0.73 1.14 0.79 1.14 0.79 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.75 0.06 0.75 0.45 0.69 0.45 0.69 0.06 0.335 0.06 0.335 0.445 0.275 0.445 0.275 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.865 0.765 0.805 0.765 0.805 0.575 0.5 0.575 0.5 1.27 0.04 1.27 0.04 1.21 0.44 1.21 0.44 0.565 0.07 0.565 0.07 0.35 0.13 0.35 0.13 0.505 0.485 0.505 0.485 0.35 0.545 0.35 0.545 0.515 0.865 0.515 ;
  END
END OR3X1

MACRO OR3X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X2 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6261 LAYER Metal1 ;
    ANTENNADIFFAREA 0.837875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.702564 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 87.923077 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.165 0.705 1.085 0.705 1.085 0.97 0.99 0.97 0.99 1.3 0.93 1.3 0.93 0.91 1.025 0.91 1.025 0.23 1.085 0.23 1.085 0.625 1.165 0.625 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.785 0.705 0.735 0.705 0.735 0.875 0.655 0.875 0.655 0.625 0.785 0.625 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.68518525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.285 0.73 0.365 1.065 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.22222225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.595 0.14 0.905 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.725 1.65 0.725 1.165 0.785 1.165 0.785 1.65 1.185 1.65 1.185 0.91 1.245 0.91 1.245 1.65 1.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 1.29 0.06 1.29 0.49 1.23 0.49 1.23 0.06 0.76 0.06 0.76 0.26 0.82 0.26 0.82 0.32 0.7 0.32 0.7 0.06 0.335 0.06 0.335 0.35 0.275 0.35 0.275 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.925 0.65 0.865 0.65 0.865 0.525 0.525 0.525 0.525 1.27 0.04 1.27 0.04 1.21 0.465 1.21 0.465 0.51 0.07 0.51 0.07 0.255 0.13 0.255 0.13 0.45 0.525 0.45 0.525 0.255 0.585 0.255 0.585 0.465 0.925 0.465 ;
  END
END OR3X2

MACRO OR3X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X4 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.98115 LAYER Metal1 ;
    ANTENNADIFFAREA 1.2471 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.3858975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 66.74358975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.565 0.73 1.49 0.73 1.49 0.97 1.375 0.97 1.375 1.46 1.315 1.46 1.315 0.97 0.965 0.97 0.965 1.46 0.905 1.46 0.905 0.91 1.43 0.91 1.43 0.49 0.945 0.49 0.945 0.25 1.005 0.25 1.005 0.43 1.37 0.43 1.37 0.23 1.43 0.23 1.43 0.42 1.49 0.42 1.49 0.6 1.565 0.6 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.4102565 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.74 0.74 1.09 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.4 1.085 0.34 1.085 0.34 1.11 0.26 1.11 0.26 0.98 0.32 0.98 0.32 0.67 0.4 0.67 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.20512825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.61 0.14 0.94 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.7 1.65 0.7 1.195 0.76 1.195 0.76 1.65 1.11 1.65 1.11 1.07 1.17 1.07 1.17 1.65 1.52 1.65 1.52 1.07 1.58 1.07 1.58 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.65 0.06 1.65 0.49 1.59 0.49 1.59 0.06 1.195 0.06 1.195 0.26 1.255 0.26 1.255 0.32 1.135 0.32 1.135 0.06 0.765 0.06 0.765 0.49 0.705 0.49 0.705 0.06 0.355 0.06 0.355 0.35 0.295 0.35 0.295 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.33 0.64 0.56 0.64 0.56 1.27 0.165 1.27 0.165 1.46 0.105 1.46 0.105 1.21 0.5 1.21 0.5 0.51 0.09 0.51 0.09 0.25 0.15 0.25 0.15 0.45 0.5 0.45 0.5 0.25 0.56 0.25 0.56 0.58 1.33 0.58 ;
  END
END OR3X4

MACRO OR3X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X6 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3545 LAYER Metal1 ;
    ANTENNADIFFAREA 2.11705 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.71794875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 59.17948725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.705 0.66 2.34 0.66 2.34 0.73 2.32 0.73 2.32 0.915 2.545 0.915 2.545 1.37 2.485 1.37 2.485 0.975 2.135 0.975 2.135 1.37 2.075 1.37 2.075 0.975 1.725 0.975 1.725 1.37 1.665 1.37 1.665 0.915 2.26 0.915 2.26 0.655 1.765 0.655 1.765 0.35 1.825 0.35 1.825 0.595 2.235 0.595 2.235 0.35 2.295 0.35 2.295 0.595 2.34 0.595 2.34 0.6 2.645 0.6 2.645 0.35 2.705 0.35 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.96 0.93 0.74 0.93 0.74 1.13 0.66 1.13 0.66 0.85 0.96 0.85 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.5897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.225 0.81 1.14 0.81 1.14 0.92 1.06 0.92 1.06 0.75 0.56 0.75 0.56 0.69 1.225 0.69 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.39 0.74 1.33 0.74 1.33 0.59 0.34 0.59 0.34 0.73 0.26 0.73 0.26 0.53 1.39 0.53 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 1.77 0 1.77 0 1.65 0.355 1.65 0.355 0.98 0.415 0.98 0.415 1.65 1.46 1.65 1.46 1.25 1.52 1.25 1.52 1.65 1.87 1.65 1.87 1.075 1.93 1.075 1.93 1.65 2.28 1.65 2.28 1.075 2.34 1.075 2.34 1.65 2.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 0.06 2.5 0.06 2.5 0.47 2.44 0.47 2.44 0.06 2.03 0.06 2.03 0.47 1.97 0.47 1.97 0.06 1.56 0.06 1.56 0.16 1.62 0.16 1.62 0.22 1.5 0.22 1.5 0.06 1.09 0.06 1.09 0.16 1.15 0.16 1.15 0.22 1.03 0.22 1.03 0.06 0.62 0.06 0.62 0.16 0.68 0.16 0.68 0.22 0.56 0.22 0.56 0.06 0.21 0.06 0.21 0.43 0.15 0.43 0.15 0.06 0 0.06 0 -0.06 2.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.1 0.815 1.55 0.815 1.55 1.09 0.99 1.09 0.99 1.37 0.93 1.37 0.93 1.03 1.49 1.03 1.49 0.43 0.325 0.43 0.325 0.37 1.55 0.37 1.55 0.755 2.1 0.755 ;
  END
END OR3X6

MACRO OR3X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3X8 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.57445 LAYER Metal1 ;
    ANTENNADIFFAREA 2.3937 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.75439725 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 51.904762 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.055 0.63 2.98 0.63 2.98 0.645 2.74 0.645 2.74 0.73 2.72 0.73 2.72 0.905 2.925 0.905 2.925 1.345 2.865 1.345 2.865 0.965 2.515 0.965 2.515 1.345 2.455 1.345 2.455 0.965 2.105 0.965 2.105 1.345 2.045 1.345 2.045 0.965 1.695 0.965 1.695 1.345 1.635 1.345 1.635 0.905 2.66 0.905 2.66 0.645 1.78 0.645 1.78 0.63 1.705 0.63 1.705 0.57 1.825 0.57 1.825 0.585 2.115 0.585 2.115 0.57 2.235 0.57 2.235 0.585 2.555 0.585 2.555 0.525 2.615 0.525 2.615 0.585 2.935 0.585 2.935 0.57 3.055 0.57 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.955 0.905 0.74 0.905 0.74 1.11 0.66 1.11 0.66 0.825 0.955 0.825 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.71794875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.195 0.785 1.14 0.785 1.14 0.92 1.06 0.92 1.06 0.725 0.53 0.725 0.53 0.665 1.195 0.665 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.76923075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.36 0.755 1.3 0.755 1.3 0.565 0.34 0.565 0.34 0.73 0.26 0.73 0.26 0.52 0.295 0.52 0.295 0.505 1.36 0.505 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 1.77 0 1.77 0 1.65 0.325 1.65 0.325 0.955 0.385 0.955 0.385 1.65 1.43 1.65 1.43 1.225 1.49 1.225 1.49 1.65 1.84 1.65 1.84 1.065 1.9 1.065 1.9 1.65 2.25 1.65 2.25 1.065 2.31 1.065 2.31 1.65 2.66 1.65 2.66 1.065 2.72 1.065 2.72 1.65 3.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 0.06 2.82 0.06 2.82 0.485 2.76 0.485 2.76 0.06 2.41 0.06 2.41 0.485 2.35 0.485 2.35 0.06 2 0.06 2 0.485 1.94 0.485 1.94 0.06 1.53 0.06 1.53 0.16 1.59 0.16 1.59 0.22 1.47 0.22 1.47 0.06 1.06 0.06 1.06 0.16 1.12 0.16 1.12 0.22 1 0.22 1 0.06 0.59 0.06 0.59 0.16 0.65 0.16 0.65 0.22 0.53 0.22 0.53 0.06 0.18 0.06 0.18 0.42 0.12 0.42 0.12 0.06 0 0.06 0 -0.06 3.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.505 0.805 1.52 0.805 1.52 1.08 0.96 1.08 0.96 1.345 0.9 1.345 0.9 1.02 1.46 1.02 1.46 0.405 0.295 0.405 0.295 0.345 1.52 0.345 1.52 0.745 2.505 0.745 ;
  END
END OR3X8

MACRO OR3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3XL 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4947 LAYER Metal1 ;
    ANTENNADIFFAREA 0.560175 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 30.537037 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 249.074074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.975 1.11 0.96 1.11 0.96 1.305 0.86 1.305 0.86 1.03 0.895 1.03 0.895 0.26 0.975 0.26 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.765 1.085 0.625 1.085 0.625 0.645 0.74 0.645 0.74 0.99 0.765 0.99 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.962963 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.64 0.405 0.925 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.462963 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.585 0.175 0.765 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.675 1.65 0.675 1.185 0.735 1.185 0.735 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.75 0.06 0.75 0.355 0.69 0.355 0.69 0.06 0.335 0.06 0.335 0.355 0.275 0.355 0.275 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.825 0.575 0.765 0.575 0.765 0.515 0.525 0.515 0.525 1.275 0.04 1.275 0.04 1.215 0.465 1.215 0.465 0.515 0.07 0.515 0.07 0.26 0.13 0.26 0.13 0.455 0.48 0.455 0.48 0.26 0.54 0.26 0.54 0.455 0.825 0.455 ;
  END
END OR3XL

MACRO OR4X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X1 0 0 ;
  SIZE 1.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.5282 LAYER Metal1 ;
    ANTENNADIFFAREA 0.73875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.05811975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 139.79487175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.155 0.54 1.115 0.54 1.115 1.385 1.055 1.385 1.055 0.275 1.115 0.275 1.115 0.41 1.155 0.41 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.55 1.07 0.5 1.07 0.5 1.11 0.42 1.11 0.42 0.98 0.47 0.98 0.47 0.66 0.55 0.66 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.62962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.37 0.87 0.3 0.87 0.3 0.96 0.22 0.96 0.22 0.79 0.29 0.79 0.29 0.59 0.37 0.59 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.9444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.16 0.705 0.15 0.705 0.15 0.84 0.09 0.84 0.09 0.705 0.08 0.705 0.08 0.545 0.16 0.545 ;
    END
  END D
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.29629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.955 0.765 0.755 0.765 0.755 0.685 0.875 0.685 0.875 0.625 0.955 0.625 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.77 0 1.77 0 1.65 0.79 1.65 0.79 1.46 0.85 1.46 0.85 1.045 0.91 1.045 0.91 1.65 1.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.06 0.91 0.06 0.91 0.495 0.85 0.495 0.85 0.06 0.56 0.06 0.56 0.2 0.44 0.2 0.44 0.06 0.17 0.06 0.17 0.2 0.04 0.2 0.04 0.06 0 0.06 0 -0.06 1.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.97 0.925 0.695 0.925 0.695 1.27 0.15 1.27 0.15 1.14 0.21 1.14 0.21 1.21 0.635 1.21 0.635 0.49 0.235 0.49 0.235 0.37 0.295 0.37 0.295 0.43 0.635 0.43 0.635 0.37 0.695 0.37 0.695 0.865 0.97 0.865 ;
  END
END OR4X1

MACRO OR4X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7968 LAYER Metal1 ;
    ANTENNADIFFAREA 1.155525 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.62051275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 103.5641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.4 1.74 1.355 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.92 0.75 0.84 0.75 0.84 0.68 0.74 0.68 0.74 0.73 0.66 0.73 0.66 0.6 0.84 0.6 0.84 0.48 0.92 0.48 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 0.96 0.46 0.96 0.46 0.79 0.48 0.79 0.48 0.48 0.56 0.48 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.36 0.96 0.26 0.96 0.26 0.79 0.28 0.79 0.28 0.48 0.36 0.48 ;
    END
  END D
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 0.705 1.275 0.705 1.275 0.76 1.195 0.76 1.195 0.35 1.275 0.35 1.275 0.625 1.365 0.625 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 1.455 1.65 1.455 1.025 1.515 1.025 1.515 1.65 1.865 1.65 1.865 0.965 1.925 0.965 1.925 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.925 0.06 1.925 0.38 1.865 0.38 1.865 0.06 1.515 0.06 1.515 0.38 1.455 0.38 1.455 0.06 0.72 0.06 0.72 0.2 0.66 0.2 0.66 0.06 0.28 0.06 0.28 0.38 0.22 0.38 0.22 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.56 0.925 1.08 0.925 1.08 1.12 0.325 1.12 0.325 1.18 0.265 1.18 0.265 1.06 1.02 1.06 1.02 0.38 0.425 0.38 0.425 0.26 0.485 0.26 0.485 0.32 1.02 0.32 1.02 0.26 1.08 0.26 1.08 0.865 1.5 0.865 1.5 0.805 1.56 0.805 ;
  END
END OR4X2

MACRO OR4X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X4 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9081 LAYER Metal1 ;
    ANTENNADIFFAREA 1.53745 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.7615385 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 62.5897435 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 1.3 1.855 1.3 1.855 1.36 1.795 1.36 1.795 1.05 1.445 1.05 1.445 1.36 1.385 1.36 1.385 0.99 1.88 0.99 1.88 0.545 1.44 0.545 1.44 0.405 1.5 0.405 1.5 0.485 1.85 0.485 1.85 0.405 1.94 0.405 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.745 0.92 0.74 0.92 0.74 1.14 0.66 1.14 0.66 0.79 0.665 0.79 0.665 0.645 0.745 0.645 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 1.125 0.46 1.125 0.46 0.8 0.48 0.8 0.48 0.645 0.56 0.645 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.61 0.34 1.11 ;
    END
  END D
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.73 1.005 0.73 1.005 0.65 1.26 0.65 1.26 0.485 1.34 0.485 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 1.11 1.65 1.11 0.99 1.17 0.99 1.17 1.65 1.59 1.65 1.59 1.24 1.65 1.24 1.65 1.65 2.04 1.65 2.04 0.97 2.1 0.97 2.1 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 2.115 0.06 2.115 0.385 2.055 0.385 2.055 0.06 1.705 0.06 1.705 0.385 1.645 0.385 1.645 0.06 1.17 0.06 1.17 0.385 1.11 0.385 1.11 0.06 0.705 0.06 0.705 0.385 0.645 0.385 0.645 0.06 0.295 0.06 0.295 0.385 0.235 0.385 0.235 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.78 0.89 0.905 0.89 0.905 1.3 0.325 1.3 0.325 1.36 0.265 1.36 0.265 1.24 0.845 1.24 0.845 0.545 0.44 0.545 0.44 0.405 0.5 0.405 0.5 0.485 0.85 0.485 0.85 0.405 0.91 0.405 0.91 0.545 0.905 0.545 0.905 0.83 1.72 0.83 1.72 0.77 1.78 0.77 ;
  END
END OR4X4

MACRO OR4X6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X6 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4884 LAYER Metal1 ;
    ANTENNADIFFAREA 2.3287 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.48091175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 62.5128205 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.97 0.585 2.72 0.585 2.72 0.98 2.74 0.98 2.74 1.05 2.88 1.05 2.88 1.37 2.82 1.37 2.82 1.11 2.47 1.11 2.47 1.37 2.41 1.37 2.41 1.04 2.06 1.04 2.06 1.37 2 1.37 2 0.98 2.66 0.98 2.66 0.585 2.09 0.585 2.09 0.275 2.15 0.275 2.15 0.525 2.5 0.525 2.5 0.275 2.56 0.275 2.56 0.525 2.91 0.525 2.91 0.275 2.97 0.275 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.74 1.11 1.72 1.11 1.72 1.23 0.3 1.23 0.3 0.89 0.36 0.89 0.36 1.17 1.66 1.17 1.66 0.805 1.72 0.805 1.72 0.98 1.74 0.98 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.69230775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.56 1.07 0.46 1.07 0.46 0.79 0.54 0.79 0.54 0.92 0.58 0.92 0.58 1.01 1.5 1.01 1.5 0.89 1.56 0.89 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 0.91 0.68 0.91 0.68 0.85 1.305 0.85 1.305 0.705 1.235 0.705 1.235 0.625 1.365 0.625 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.135 0.75 0.68 0.75 0.68 0.625 0.965 0.625 0.965 0.67 1.135 0.67 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 1.77 0 1.77 0 1.65 0.255 1.65 0.255 1.33 0.315 1.33 0.315 1.65 1.735 1.65 1.735 1.54 1.855 1.54 1.855 1.65 2.205 1.65 2.205 1.14 2.265 1.14 2.265 1.65 2.615 1.65 2.615 1.21 2.675 1.21 2.675 1.65 3.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 0.06 2.765 0.06 2.765 0.395 2.705 0.395 2.705 0.06 2.355 0.06 2.355 0.395 2.295 0.395 2.295 0.06 1.915 0.06 1.915 0.305 1.975 0.305 1.975 0.365 1.855 0.365 1.855 0.06 1.475 0.06 1.475 0.305 1.535 0.305 1.535 0.365 1.415 0.365 1.415 0.06 1.035 0.06 1.035 0.305 1.095 0.305 1.095 0.365 0.975 0.365 0.975 0.06 0.595 0.06 0.595 0.305 0.655 0.305 0.655 0.365 0.535 0.365 0.535 0.06 0.2 0.06 0.2 0.395 0.14 0.395 0.14 0.06 0 0.06 0 -0.06 3.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.425 0.75 1.9 0.75 1.9 1.39 1.04 1.39 1.04 1.33 1.84 1.33 1.84 0.525 0.385 0.525 0.385 0.505 0.315 0.505 0.315 0.445 0.435 0.445 0.435 0.465 0.755 0.465 0.755 0.445 0.875 0.445 0.875 0.465 1.195 0.465 1.195 0.445 1.315 0.445 1.315 0.465 1.635 0.465 1.635 0.445 1.755 0.445 1.755 0.465 1.9 0.465 1.9 0.69 2.425 0.69 ;
  END
END OR4X6

MACRO OR4X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4X8 0 0 ;
  SIZE 3.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.74155 LAYER Metal1 ;
    ANTENNADIFFAREA 2.636775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2331 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.471257 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 56.3835265 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.41 0.54 3.335 0.54 3.335 0.555 3.14 0.555 3.14 0.815 3.315 0.815 3.315 1.345 3.255 1.345 3.255 0.875 2.905 0.875 2.905 1.345 2.845 1.345 2.845 0.875 2.495 0.875 2.495 1.345 2.435 1.345 2.435 0.875 2.085 0.875 2.085 1.345 2.025 1.345 2.025 0.815 3.06 0.815 3.06 0.555 2.135 0.555 2.135 0.54 2.06 0.54 2.06 0.48 2.18 0.48 2.18 0.495 2.47 0.495 2.47 0.48 2.59 0.48 2.59 0.495 2.91 0.495 2.91 0.435 2.97 0.435 2.97 0.495 3.29 0.495 3.29 0.48 3.41 0.48 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.5641025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.765 0.895 1.695 0.895 1.695 1.23 0.27 1.23 0.27 0.865 0.33 0.865 0.33 1.17 1.635 1.17 1.635 0.775 1.74 0.775 1.74 0.815 1.765 0.815 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5128205 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.535 1.07 0.46 1.07 0.46 0.79 0.54 0.79 0.54 0.92 0.58 0.92 0.58 1.01 1.475 1.01 1.475 0.9 1.535 0.9 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 0.91 0.68 0.91 0.68 0.85 1.305 0.85 1.305 0.705 1.235 0.705 1.235 0.625 1.365 0.625 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.974359 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.135 0.75 0.68 0.75 0.68 0.625 0.965 0.625 0.965 0.67 1.135 0.67 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 1.77 0 1.77 0 1.65 0.255 1.65 0.255 1.33 0.315 1.33 0.315 1.65 1.755 1.65 1.755 1.54 1.875 1.54 1.875 1.65 2.23 1.65 2.23 0.975 2.29 0.975 2.29 1.65 2.64 1.65 2.64 0.975 2.7 0.975 2.7 1.65 3.05 1.65 3.05 1.065 3.11 1.065 3.11 1.65 3.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 0.06 3.175 0.06 3.175 0.395 3.115 0.395 3.115 0.06 2.765 0.06 2.765 0.395 2.705 0.395 2.705 0.06 2.355 0.06 2.355 0.395 2.295 0.395 2.295 0.06 1.915 0.06 1.915 0.305 1.975 0.305 1.975 0.365 1.855 0.365 1.855 0.06 1.475 0.06 1.475 0.305 1.535 0.305 1.535 0.365 1.415 0.365 1.415 0.06 1.035 0.06 1.035 0.305 1.095 0.305 1.095 0.365 0.975 0.365 0.975 0.06 0.595 0.06 0.595 0.305 0.655 0.305 0.655 0.365 0.535 0.365 0.535 0.06 0.2 0.06 0.2 0.395 0.14 0.395 0.14 0.06 0 0.06 0 -0.06 3.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.86 0.715 1.925 0.715 1.925 1.39 1.04 1.39 1.04 1.33 1.865 1.33 1.865 0.525 0.385 0.525 0.385 0.505 0.315 0.505 0.315 0.445 0.435 0.445 0.435 0.465 0.755 0.465 0.755 0.445 0.875 0.445 0.875 0.465 1.195 0.465 1.195 0.445 1.315 0.445 1.315 0.465 1.635 0.465 1.635 0.445 1.755 0.445 1.755 0.465 1.925 0.465 1.925 0.655 2.86 0.655 ;
  END
END OR4X8

MACRO OR4XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR4XL 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6027 LAYER Metal1 ;
    ANTENNADIFFAREA 0.827725 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXAREACAR 37.20370375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 283.611111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.37 1.54 1.315 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.755 1.085 0.675 1.085 0.675 0.73 0.66 0.73 0.66 0.6 0.74 0.6 0.74 0.65 0.755 0.65 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.56 1.11 0.46 1.11 0.46 0.98 0.48 0.98 0.48 0.63 0.56 0.63 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.6 0.34 1.1 ;
    END
  END D
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 1.03 1.12 1.03 1.12 0.73 1.06 0.73 1.06 0.59 1.2 0.59 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 1.135 1.65 1.135 1.29 1.195 1.29 1.195 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.25 0.06 1.25 0.49 1.19 0.49 1.19 0.06 0.72 0.06 0.72 0.2 0.66 0.2 0.66 0.06 0.32 0.06 0.32 0.2 0.26 0.2 0.26 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.36 1.19 0.915 1.19 0.915 1.285 0.235 1.285 0.235 1.225 0.855 1.225 0.855 0.49 0.425 0.49 0.425 0.37 0.485 0.37 0.485 0.43 0.855 0.43 0.855 0.37 0.915 0.37 0.915 1.13 1.3 1.13 1.3 1.025 1.36 1.025 ;
  END
END OR4XL

MACRO PBUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN PBUFX2 0 0 ;
  SIZE 2.8 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.04 2.445 1.98 2.445 1.98 1.94 1.63 1.94 1.63 2.445 1.57 2.445 1.57 1.94 1.405 1.94 1.405 2.63 0.955 2.63 0.955 2.035 1.015 2.035 1.015 2.31 1.345 2.31 1.345 1.88 2.04 1.88 ;
    END
  END ExtVDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.405 2.485 0.64 2.655 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8172 LAYER Metal1 ;
    ANTENNADIFFAREA 0.766 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.96923075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 103.076923 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.03 2.82 1.835 2.82 1.835 3.16 1.775 3.16 1.775 2.055 1.835 2.055 1.835 2.69 2.03 2.69 ;
    END
  END Y
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 3.48 0 3.48 0 3.36 0.955 3.36 0.955 2.97 1.015 2.97 1.015 3.36 1.57 3.36 1.57 2.9 1.63 2.9 1.63 3.36 1.98 3.36 1.98 2.9 2.04 2.9 2.04 3.36 2.8 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 2.8 0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 2.8 1.77 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.69 2.79 0.81 2.79 0.81 3.115 0.75 3.115 0.75 2.035 0.81 2.035 0.81 2.73 1.69 2.73 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
  PROPERTY vceLastSavedModifiedCounter 8926 ;
END PBUFX2

MACRO PINVX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN PINVX1 0 0 ;
  SIZE 2.2 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.4568 LAYER Metal1 ;
    ANTENNADIFFAREA 0.5006 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.87 1.94 0.93 3.15 ;
    END
  END Y
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.625 2.63 1.075 2.63 1.075 1.94 1.275 1.94 1.275 2.33 1.135 2.33 1.135 2.49 1.625 2.49 ;
    END
  END ExtVDD
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.56 2.69 0.745 2.82 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 3.48 0 3.48 0 3.36 1.075 3.36 1.075 2.89 1.135 2.89 1.135 3.36 2.2 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        RECT 0 -0.06 2.2 0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 0 1.65 2.2 1.77 ;
    END
  END VDD
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END PINVX1

MACRO RDFFNQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RDFFNQX1 0 0 ;
  SIZE 4.6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.77 4.365 1.77 4.365 2.46 4.305 2.46 4.305 1.77 1.035 1.77 1.035 2.4 0.975 2.4 0.975 1.77 0.255 1.77 0.255 2.4 0.195 2.4 0.195 1.77 0 1.77 0 1.65 0.895 1.65 0.895 1.11 0.955 1.11 0.955 1.65 4.3 1.65 4.3 1.13 4.36 1.13 4.36 1.65 4.6 1.65 ;
    END
  END VDD
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.9 2.61 2.42 2.61 2.42 2 2.57 2 2.57 1.89 2.82 1.89 2.82 2 2.9 2 ;
    END
  END ExtVDD
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8127 LAYER Metal1 ;
    ANTENNADIFFAREA 2.739875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20745 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.3788865 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 132.8850325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.165 2.83 4.16 2.83 4.16 3.135 4.1 3.135 4.1 2.83 4.03 2.83 4.03 2.68 4.1 2.68 4.1 2.07 4.16 2.07 4.16 2.68 4.165 2.68 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.87037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.11 2.46 0.365 2.63 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 3.48 0 3.48 0 3.36 0.195 3.36 0.195 2.97 0.255 2.97 0.255 3.36 0.975 3.36 0.975 2.97 1.035 2.97 1.035 3.36 2.42 3.36 2.42 3.025 2.48 3.025 2.48 3.36 2.84 3.36 2.84 3.025 2.9 3.025 2.9 3.36 4.305 3.36 4.305 2.875 4.365 2.875 4.365 3.36 4.6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 0.06 4.36 0.06 4.36 0.465 4.3 0.465 4.3 0.06 2.995 0.06 2.995 0.625 2.935 0.625 2.935 0.06 0.955 0.06 0.955 0.54 0.895 0.54 0.895 0.06 0 0.06 0 -0.06 4.6 -0.06 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.9444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.935 2.5 1.165 2.645 ;
    END
  END CKN
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0993 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 3.06481475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 23.425926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.46 1.13 3.7 1.36 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 4.05 1.345 3.99 1.345 3.99 1.05 3.96 1.05 3.96 0.93 3.99 0.93 3.99 0.32 4.05 0.32 ;
      RECT 3.775 0.14 3.835 1.45 ;
      RECT 3.3 2.615 3.745 2.675 ;
      POLYGON 3.42 1.525 3.14 1.525 3.14 1.025 2.66 1.025 2.66 0.38 2.72 0.38 2.72 0.965 3.14 0.965 3.14 0.48 3.2 0.48 3.2 1.465 3.42 1.465 ;
      RECT 3.31 0.48 3.37 1.215 ;
      POLYGON 3.21 3.17 3.15 3.17 3.15 2.78 2.35 2.78 2.35 2.72 3.15 2.72 3.15 2 3.21 2 ;
      POLYGON 3.005 2.93 2.275 2.93 2.275 3.17 2.215 3.17 2.215 2 2.275 2 2.275 2.87 3.005 2.87 ;
      POLYGON 2.995 1.555 2.735 1.555 2.735 1.26 2.935 1.26 2.935 1.255 2.995 1.255 ;
      RECT 2.42 0.48 2.48 1.47 ;
      POLYGON 2.275 1.54 2.005 1.54 2.005 1.48 2.215 1.48 2.215 0.48 2.275 0.48 ;
      POLYGON 2.125 1.02 2.005 1.02 2.005 0.96 2.035 0.96 2.035 0.86 1.365 0.86 1.365 1.325 1.305 1.325 1.305 0.38 1.365 0.38 1.365 0.8 2.095 0.8 2.095 0.96 2.125 0.96 ;
      POLYGON 1.3 3.03 1.24 3.03 1.24 3.115 1.18 3.115 1.18 2.97 1.24 2.97 1.24 2.795 0.895 2.795 0.895 2.735 1.24 2.735 1.24 2.4 1.18 2.4 1.18 2.185 1.24 2.185 1.24 2.25 1.3 2.25 ;
      POLYGON 1.16 1.325 1.1 1.325 1.1 0.85 0.89 0.85 0.89 0.98 0.92 0.98 0.92 1.04 0.8 1.04 0.8 0.98 0.83 0.98 0.83 0.67 0.8 0.67 0.8 0.61 0.92 0.61 0.92 0.67 0.89 0.67 0.89 0.79 1.1 0.79 1.1 0.395 1.16 0.395 ;
      POLYGON 0.83 3.115 0.77 3.115 0.77 2.795 0.68 2.795 0.68 2.735 0.77 2.735 0.77 1.885 0.83 1.885 ;
      POLYGON 0.645 1.325 0.635 1.325 0.635 1.525 0.475 1.525 0.475 1.465 0.575 1.465 0.575 1.11 0.585 1.11 0.585 0.395 0.645 0.395 ;
      POLYGON 0.61 2.155 0.565 2.155 0.565 3.115 0.505 3.115 0.505 2.095 0.55 2.095 0.55 1.84 0.61 1.84 ;
      RECT 0.305 0.145 0.365 1.545 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RDFFNQX1

MACRO RDFFNRQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RDFFNRQX1 0 0 ;
  SIZE 5.6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 5.185 1.77 5.185 2.46 5.125 2.46 5.125 1.77 1.56 1.77 1.56 2.385 1.5 2.385 1.5 1.77 1.115 1.77 1.115 2.4 1.055 2.4 1.055 1.77 0.26 1.77 0.26 2.4 0.2 2.4 0.2 1.77 -0.005 1.77 -0.005 1.65 0.89 1.65 0.89 1.27 0.95 1.27 0.95 1.65 1.44 1.65 1.44 1.27 1.5 1.27 1.5 1.65 5.03 1.65 5.03 1.13 5.09 1.13 5.09 1.65 5.6 1.65 ;
    END
  END VDD
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.495 2.61 3.015 2.61 3.015 2 3.145 2 3.145 1.89 3.395 1.89 3.395 2 3.495 2 ;
    END
  END ExtVDD
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.03 2.69 1.185 2.845 ;
    END
  END CKN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.31481475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.64 2.59 1.63 2.59 1.63 2.655 1.415 2.655 1.415 2.485 1.63 2.485 1.63 2.53 1.64 2.53 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.54205 LAYER Metal1 ;
    ANTENNADIFFAREA 3.382925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.23985 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.937044 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 138.4615385 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.98 3.135 4.92 3.135 4.92 2.765 4.835 2.765 4.835 2.635 4.92 2.635 4.92 2.07 4.98 2.07 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.16 2.5 0.355 2.63 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 3.48 0 3.48 0 3.36 0.2 3.36 0.2 2.97 0.26 2.97 0.26 3.36 1.055 3.36 1.055 2.97 1.115 2.97 1.115 3.36 1.5 3.36 1.5 2.97 1.56 2.97 1.56 3.36 3.015 3.36 3.015 3.025 3.075 3.025 3.075 3.36 3.435 3.36 3.435 3.025 3.495 3.025 3.495 3.36 5.125 3.36 5.125 2.875 5.185 2.875 5.185 3.36 5.6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5.46 0.06 5.46 0.465 5.4 0.465 5.4 0.06 5.05 0.06 5.05 0.465 4.99 0.465 4.99 0.06 3.59 0.06 3.59 0.465 3.53 0.465 3.53 0.06 1.405 0.06 1.405 0.465 1.345 0.465 1.345 0.06 0.95 0.06 0.95 0.465 0.89 0.465 0.89 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.10185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.21 1.525 4.055 1.525 4.055 1.37 3.91 1.37 3.91 0.41 3.97 0.41 3.97 1.31 4.21 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.4 1.345 5.34 1.345 5.34 1.015 4.85 1.015 4.85 1.345 4.79 1.345 4.79 0.955 5.4 0.955 ;
      POLYGON 5.255 0.67 4.79 0.67 4.79 0.32 4.85 0.32 4.85 0.61 5.195 0.61 5.195 0.32 5.255 0.32 ;
      RECT 4.585 0.32 4.645 1.345 ;
      RECT 3.895 2.385 4.34 2.445 ;
      POLYGON 4.335 1.08 4.065 1.08 4.065 0.25 4.055 0.25 4.055 0.23 4.04 0.23 4.04 0.17 4.055 0.17 4.055 0.13 4.115 0.13 4.115 0.17 4.125 0.17 4.125 1.02 4.335 1.02 ;
      POLYGON 3.995 1.51 3.735 1.51 3.735 0.685 3.2 0.685 3.2 0.52 3.26 0.52 3.26 0.625 3.735 0.625 3.735 0.32 3.795 0.32 3.795 1.45 3.995 1.45 ;
      POLYGON 3.805 3.17 3.745 3.17 3.745 2.78 2.945 2.78 2.945 2.72 3.745 2.72 3.745 2 3.805 2 ;
      POLYGON 3.6 2.93 2.87 2.93 2.87 3.17 2.81 3.17 2.81 2 2.87 2 2.87 2.87 3.6 2.87 ;
      RECT 3.31 1.24 3.59 1.525 ;
      RECT 3.015 0.32 3.075 1.455 ;
      POLYGON 2.87 1.52 2.58 1.52 2.58 1.46 2.81 1.46 2.81 0.32 2.87 0.32 ;
      RECT 2.275 0.71 2.335 1.285 ;
      POLYGON 1.945 1.485 1.885 1.485 1.885 0.85 1.755 0.85 1.755 0.32 1.815 0.32 1.815 0.79 1.945 0.79 ;
      POLYGON 1.805 2.57 1.765 2.57 1.765 3.115 1.705 3.115 1.705 2.17 1.765 2.17 1.765 2.45 1.805 2.45 ;
      POLYGON 1.74 1.485 1.68 1.485 1.68 1.2 1.19 1.2 1.19 1.485 1.13 1.485 1.13 1.2 0.795 1.2 0.795 1.14 1.28 1.14 1.28 0.595 0.795 0.595 0.795 0.535 1.095 0.535 1.095 0.32 1.155 0.32 1.155 0.535 1.55 0.535 1.55 0.32 1.61 0.32 1.61 0.595 1.34 0.595 1.34 1.14 1.74 1.14 ;
      POLYGON 1.32 3.115 1.26 3.115 1.26 2.6 0.98 2.6 0.98 2.54 1.26 2.54 1.26 2.185 1.32 2.185 ;
      POLYGON 0.91 3.115 0.85 3.115 0.85 2.82 0.79 2.82 0.79 2.7 0.85 2.7 0.85 1.86 0.91 1.86 ;
      POLYGON 0.64 1.525 0.37 1.525 0.37 1.465 0.58 1.465 0.58 0.32 0.64 0.32 ;
      POLYGON 0.64 2.075 0.57 2.075 0.57 3.115 0.51 3.115 0.51 2.015 0.64 2.015 ;
      RECT 0.28 0.135 0.34 1.305 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RDFFNRQX1

MACRO RDFFNRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RDFFNRX1 0 0 ;
  SIZE 5.8 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 1.77 5.53 1.77 5.53 2.46 5.47 2.46 5.47 1.77 4.85 1.77 4.85 2.46 4.79 2.46 4.79 1.77 1.56 1.77 1.56 2.385 1.5 2.385 1.5 1.77 1.115 1.77 1.115 2.4 1.055 2.4 1.055 1.77 0.26 1.77 0.26 2.4 0.2 2.4 0.2 1.77 -0.005 1.77 -0.005 1.65 0.89 1.65 0.89 1.27 0.95 1.27 0.95 1.65 1.44 1.65 1.44 1.27 1.5 1.27 1.5 1.65 5.03 1.65 5.03 1.13 5.09 1.13 5.09 1.65 5.8 1.65 ;
    END
  END VDD
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.495 2.61 3.015 2.61 3.015 2 3.145 2 3.145 1.89 3.395 1.89 3.395 2 3.495 2 ;
    END
  END ExtVDD
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.985 2.69 1.185 2.845 ;
    END
  END CKN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.62 2.59 1.595 2.59 1.595 2.85 1.425 2.85 1.425 2.455 1.595 2.455 1.595 2.53 1.62 2.53 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8422 LAYER Metal1 ;
    ANTENNADIFFAREA 3.681325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2853 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.97230975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 125.488959 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.365 2.835 5.325 2.835 5.325 3.135 5.265 3.135 5.265 2.835 5.225 2.835 5.225 2.68 5.265 2.68 5.265 2.07 5.325 2.07 5.325 2.68 5.365 2.68 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.8422 LAYER Metal1 ;
    ANTENNADIFFAREA 3.681325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2853 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.97230975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 125.488959 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.645 3.135 4.585 3.135 4.585 2.63 4.435 2.63 4.435 2.5 4.585 2.5 4.585 2.07 4.645 2.07 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.16 2.5 0.365 2.63 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 3.48 0 3.48 0 3.36 0.2 3.36 0.2 2.97 0.26 2.97 0.26 3.36 1.055 3.36 1.055 2.97 1.115 2.97 1.115 3.36 1.5 3.36 1.5 2.97 1.56 2.97 1.56 3.36 3.015 3.36 3.015 3.025 3.075 3.025 3.075 3.36 3.435 3.36 3.435 3.025 3.495 3.025 3.495 3.36 4.79 3.36 4.79 2.875 4.85 2.875 4.85 3.36 5.47 3.36 5.47 2.875 5.53 2.875 5.53 3.36 5.8 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 0.06 5.46 0.06 5.46 0.465 5.4 0.465 5.4 0.06 5.05 0.06 5.05 0.465 4.99 0.465 4.99 0.06 3.59 0.06 3.59 0.465 3.53 0.465 3.53 0.06 1.405 0.06 1.405 0.465 1.345 0.465 1.345 0.06 0.95 0.06 0.95 0.465 0.89 0.465 0.89 0.06 0 0.06 0 -0.06 5.8 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.10185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.21 1.525 4.055 1.525 4.055 1.37 3.91 1.37 3.91 0.41 3.97 0.41 3.97 1.31 4.21 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.4 1.345 5.34 1.345 5.34 1.015 4.85 1.015 4.85 1.345 4.79 1.345 4.79 0.955 5.4 0.955 ;
      POLYGON 5.255 0.67 4.79 0.67 4.79 0.32 4.85 0.32 4.85 0.61 5.195 0.61 5.195 0.32 5.255 0.32 ;
      POLYGON 5.085 3.075 5.025 3.075 5.025 2.68 4.73 2.68 4.73 2.62 5.025 2.62 5.025 2.155 5.085 2.155 ;
      RECT 4.585 0.32 4.645 1.345 ;
      RECT 3.895 2.385 4.34 2.445 ;
      POLYGON 4.335 1.08 4.065 1.08 4.065 0.25 4.055 0.25 4.055 0.23 4.04 0.23 4.04 0.17 4.055 0.17 4.055 0.13 4.115 0.13 4.115 0.17 4.125 0.17 4.125 1.02 4.335 1.02 ;
      POLYGON 3.995 1.51 3.735 1.51 3.735 0.685 3.2 0.685 3.2 0.52 3.26 0.52 3.26 0.625 3.735 0.625 3.735 0.32 3.795 0.32 3.795 1.45 3.995 1.45 ;
      POLYGON 3.805 3.17 3.745 3.17 3.745 2.78 2.945 2.78 2.945 2.72 3.745 2.72 3.745 2 3.805 2 ;
      POLYGON 3.6 2.93 2.87 2.93 2.87 3.17 2.81 3.17 2.81 2 2.87 2 2.87 2.87 3.6 2.87 ;
      RECT 3.31 1.24 3.59 1.525 ;
      RECT 3.015 0.32 3.075 1.455 ;
      POLYGON 2.87 1.52 2.58 1.52 2.58 1.46 2.81 1.46 2.81 0.32 2.87 0.32 ;
      RECT 2.275 0.71 2.335 1.285 ;
      POLYGON 1.945 1.485 1.885 1.485 1.885 0.85 1.755 0.85 1.755 0.32 1.815 0.32 1.815 0.79 1.945 0.79 ;
      POLYGON 1.805 2.57 1.765 2.57 1.765 3.115 1.705 3.115 1.705 2.17 1.765 2.17 1.765 2.45 1.805 2.45 ;
      POLYGON 1.74 1.485 1.68 1.485 1.68 1.2 1.19 1.2 1.19 1.485 1.13 1.485 1.13 1.2 0.795 1.2 0.795 1.14 1.28 1.14 1.28 0.595 0.795 0.595 0.795 0.535 1.095 0.535 1.095 0.32 1.155 0.32 1.155 0.535 1.55 0.535 1.55 0.32 1.61 0.32 1.61 0.595 1.34 0.595 1.34 1.14 1.74 1.14 ;
      POLYGON 1.32 3.115 1.26 3.115 1.26 2.6 0.98 2.6 0.98 2.54 1.26 2.54 1.26 2.185 1.32 2.185 ;
      POLYGON 0.91 3.115 0.85 3.115 0.85 2.82 0.79 2.82 0.79 2.7 0.85 2.7 0.85 1.86 0.91 1.86 ;
      POLYGON 0.64 1.525 0.37 1.525 0.37 1.465 0.58 1.465 0.58 0.32 0.64 0.32 ;
      POLYGON 0.64 2.075 0.57 2.075 0.57 3.115 0.51 3.115 0.51 2.015 0.64 2.015 ;
      RECT 0.28 0.135 0.34 1.305 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RDFFNRX1

MACRO RDFFNSQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RDFFNSQX1 0 0 ;
  SIZE 5.6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 5.425 1.77 5.425 2.46 5.365 2.46 5.365 1.77 1.115 1.77 1.115 2.4 1.055 2.4 1.055 1.77 0.26 1.77 0.26 2.4 0.2 2.4 0.2 1.77 -0.005 1.77 -0.005 1.65 0.7 1.65 0.7 1.165 0.76 1.165 0.76 1.65 1.38 1.65 1.38 1.25 1.385 1.25 1.385 1.165 1.445 1.165 1.445 1.38 1.44 1.38 1.44 1.65 5.03 1.65 5.03 1.13 5.09 1.13 5.09 1.65 5.44 1.65 5.44 1.13 5.5 1.13 5.5 1.65 5.6 1.65 ;
    END
  END VDD
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0516 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.5925925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 22.2685185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.965 0.92 0.9 0.92 0.9 1.035 0.93 1.035 0.93 1.095 0.81 1.095 0.81 1.035 0.84 1.035 0.84 0.92 0.835 0.92 0.835 0.72 0.965 0.72 ;
    END
  END SN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.495 2.61 3.015 2.61 3.015 2 3.145 2 3.145 1.89 3.395 1.89 3.395 2 3.495 2 ;
    END
  END ExtVDD
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.03 2.69 1.185 2.845 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.55755 LAYER Metal1 ;
    ANTENNADIFFAREA 3.3359 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20745 LAYER Metal1 ;
      ANTENNAMAXAREACAR 21.96939025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 156.8185105 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.22 3.135 5.16 3.135 5.16 2.82 5.035 2.82 5.035 2.5 5.16 2.5 5.16 2.07 5.22 2.07 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.2 2.69 0.36 2.82 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 3.48 0 3.48 0 3.36 0.2 3.36 0.2 2.97 0.26 2.97 0.26 3.36 1.055 3.36 1.055 2.97 1.115 2.97 1.115 3.36 3.015 3.36 3.015 3.025 3.075 3.025 3.075 3.36 3.435 3.36 3.435 3.025 3.495 3.025 3.495 3.36 5.365 3.36 5.365 2.875 5.425 2.875 5.425 3.36 5.6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5.5 0.06 5.5 0.465 5.44 0.465 5.44 0.06 3.59 0.06 3.59 0.465 3.53 0.465 3.53 0.06 0.76 0.06 0.76 0.32 0.935 0.32 0.935 0.465 0.7 0.465 0.7 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.10185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.21 1.525 4.055 1.525 4.055 1.37 3.91 1.37 3.91 0.41 3.97 0.41 3.97 1.31 4.21 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.295 1.345 5.235 1.345 5.235 1.015 4.85 1.015 4.85 1.345 4.79 1.345 4.79 0.955 5.295 0.955 ;
      POLYGON 5.19 0.465 5.13 0.465 5.13 0.42 4.85 0.42 4.85 0.495 4.79 0.495 4.79 0.32 4.85 0.32 4.85 0.36 5.13 0.36 5.13 0.32 5.19 0.32 ;
      RECT 4.585 0.32 4.645 1.345 ;
      RECT 3.895 2.385 4.34 2.445 ;
      POLYGON 4.335 1.13 4.065 1.13 4.065 0.25 4.055 0.25 4.055 0.23 4.04 0.23 4.04 0.17 4.055 0.17 4.055 0.13 4.115 0.13 4.115 0.17 4.125 0.17 4.125 1.07 4.335 1.07 ;
      RECT 4.245 0.135 4.305 0.995 ;
      POLYGON 3.995 1.51 3.735 1.51 3.735 0.83 3.2 0.83 3.2 0.245 3.26 0.245 3.26 0.77 3.735 0.77 3.735 0.32 3.795 0.32 3.795 1.45 3.995 1.45 ;
      POLYGON 3.805 3.17 3.745 3.17 3.745 2.78 2.945 2.78 2.945 2.72 3.745 2.72 3.745 2 3.805 2 ;
      POLYGON 3.6 2.93 2.87 2.93 2.87 3.17 2.81 3.17 2.81 2 2.87 2 2.87 2.87 3.6 2.87 ;
      RECT 3.31 1.24 3.59 1.525 ;
      RECT 3.015 0.32 3.075 1.455 ;
      POLYGON 2.87 1.52 2.58 1.52 2.58 1.46 2.81 1.46 2.81 0.32 2.87 0.32 ;
      RECT 2.275 0.6 2.335 1.18 ;
      POLYGON 1.95 0.83 1.89 0.83 1.89 1.38 1.83 1.38 1.83 0.32 1.89 0.32 1.89 0.77 1.95 0.77 ;
      POLYGON 1.685 1.38 1.625 1.38 1.625 0.585 1.12 0.585 1.12 1.165 1.24 1.165 1.24 1.38 0.905 1.38 0.905 1.165 1.06 1.165 1.06 0.585 0.725 0.585 0.725 0.595 0.695 0.595 0.695 1.035 0.725 1.035 0.725 1.095 0.605 1.095 0.605 1.035 0.635 1.035 0.635 0.595 0.605 0.595 0.605 0.535 0.635 0.535 0.635 0.525 1.185 0.525 1.185 0.32 1.245 0.32 1.245 0.525 1.625 0.525 1.625 0.32 1.685 0.32 ;
      POLYGON 1.335 0.705 1.305 0.705 1.305 1.035 1.335 1.035 1.335 1.095 1.215 1.095 1.215 1.035 1.245 1.035 1.245 0.705 1.215 0.705 1.215 0.645 1.335 0.645 ;
      POLYGON 1.32 3.115 1.26 3.115 1.26 2.6 0.98 2.6 0.98 2.54 1.26 2.54 1.26 2.185 1.32 2.185 ;
      POLYGON 0.91 3.115 0.85 3.115 0.85 2.82 0.79 2.82 0.79 2.7 0.85 2.7 0.85 1.86 0.91 1.86 ;
      POLYGON 0.64 2.1 0.57 2.1 0.57 3.115 0.51 3.115 0.51 2.015 0.61 2.015 0.61 2.04 0.64 2.04 ;
      POLYGON 0.45 1.52 0.29 1.52 0.29 1.46 0.39 1.46 0.39 0.32 0.45 0.32 ;
      RECT 0.1 0.135 0.16 1.2 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RDFFNSQX1

MACRO RDFFNSRQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RDFFNSRQX1 0 0 ;
  SIZE 6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 1.77 5.73 1.77 5.73 2.46 5.67 2.46 5.67 1.77 1.56 1.77 1.56 2.385 1.5 2.385 1.5 1.77 1.115 1.77 1.115 2.4 1.055 2.4 1.055 1.77 0.26 1.77 0.26 2.4 0.2 2.4 0.2 1.77 -0.005 1.77 -0.005 1.65 0.89 1.65 0.89 1.27 0.95 1.27 0.95 1.65 1.68 1.65 1.68 1.27 1.74 1.27 1.74 1.65 5.23 1.65 5.23 1.13 5.29 1.13 5.29 1.65 5.745 1.65 5.745 1.13 5.805 1.13 5.805 1.65 6 1.65 ;
    END
  END VDD
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0516 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.5925925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 23.287037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.165 0.92 1.09 0.92 1.09 1.14 1.12 1.14 1.12 1.2 1 1.2 1 1.14 1.03 1.14 1.03 0.72 1.165 0.72 ;
    END
  END SN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.695 2.61 3.215 2.61 3.215 2 3.345 2 3.345 1.89 3.595 1.89 3.595 2 3.695 2 ;
    END
  END ExtVDD
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.64814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 2.69 1.185 2.845 ;
    END
  END CKN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.64814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 2.5 1.61 2.63 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.047325 LAYER Metal1 ;
    ANTENNADIFFAREA 3.6339 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.23985 LAYER Metal1 ;
      ANTENNAMAXAREACAR 21.04367325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 154.15884925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.565 2.82 5.525 2.82 5.525 3.135 5.465 3.135 5.465 2.82 5.435 2.82 5.435 2.5 5.465 2.5 5.465 2.07 5.525 2.07 5.525 2.5 5.565 2.5 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.462963 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.2 2.495 0.365 2.625 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 3.48 0 3.48 0 3.36 0.2 3.36 0.2 2.97 0.26 2.97 0.26 3.36 1.055 3.36 1.055 2.97 1.115 2.97 1.115 3.36 1.5 3.36 1.5 2.97 1.56 2.97 1.56 3.36 3.215 3.36 3.215 3.025 3.275 3.025 3.275 3.36 3.635 3.36 3.635 3.025 3.695 3.025 3.695 3.36 5.67 3.36 5.67 2.875 5.73 2.875 5.73 3.36 6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6 0.06 5.865 0.06 5.865 0.465 5.805 0.465 5.805 0.06 3.79 0.06 3.79 0.465 3.73 0.465 3.73 0.06 0.95 0.06 0.95 0.32 1.125 0.32 1.125 0.465 0.89 0.465 0.89 0.06 0 0.06 0 -0.06 6 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.537037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.565 1.525 4.275 1.525 4.275 1.36 4.11 1.36 4.11 0.41 4.17 0.41 4.17 1.3 4.335 1.3 4.335 1.36 4.565 1.36 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.66 0.465 5.6 0.465 5.6 0.26 5.25 0.26 5.25 0.465 5.19 0.465 5.19 0.2 5.66 0.2 ;
      POLYGON 5.6 1.345 5.54 1.345 5.54 1.015 5.05 1.015 5.05 1.345 4.99 1.345 4.99 0.955 5.6 0.955 ;
      POLYGON 5.455 0.67 4.99 0.67 4.99 0.32 5.05 0.32 5.05 0.61 5.395 0.61 5.395 0.32 5.455 0.32 ;
      RECT 4.785 0.32 4.845 1.345 ;
      RECT 4.095 2.385 4.54 2.445 ;
      POLYGON 4.535 1.13 4.265 1.13 4.265 0.25 4.255 0.25 4.255 0.23 4.24 0.23 4.24 0.17 4.255 0.17 4.255 0.13 4.315 0.13 4.315 0.17 4.325 0.17 4.325 1.07 4.535 1.07 ;
      RECT 4.445 0.135 4.505 0.995 ;
      POLYGON 4.205 1.51 3.935 1.51 3.935 0.83 3.4 0.83 3.4 0.245 3.46 0.245 3.46 0.77 3.935 0.77 3.935 0.32 3.995 0.32 3.995 1.45 4.205 1.45 ;
      POLYGON 4.005 3.17 3.945 3.17 3.945 2.78 3.145 2.78 3.145 2.72 3.945 2.72 3.945 2 4.005 2 ;
      POLYGON 3.8 2.93 3.07 2.93 3.07 3.17 3.01 3.17 3.01 2 3.07 2 3.07 2.87 3.8 2.87 ;
      RECT 3.51 1.24 3.79 1.525 ;
      RECT 3.215 0.32 3.275 1.455 ;
      POLYGON 3.07 1.52 2.78 1.52 2.78 1.46 3.01 1.46 3.01 0.32 3.07 0.32 ;
      RECT 2.475 0.6 2.535 1.285 ;
      POLYGON 2.245 0.83 2.185 0.83 2.185 1.485 2.125 1.485 2.125 0.32 2.185 0.32 2.185 0.77 2.245 0.77 ;
      POLYGON 2.065 1.19 1.98 1.19 1.98 1.485 1.92 1.485 1.92 1.13 2.005 1.13 2.005 0.585 1.31 0.585 1.31 1.27 1.43 1.27 1.43 1.485 1.095 1.485 1.095 1.27 1.25 1.27 1.25 0.585 0.915 0.585 0.915 0.595 0.885 0.595 0.885 1.14 0.915 1.14 0.915 1.2 0.795 1.2 0.795 1.14 0.825 1.14 0.825 0.595 0.795 0.595 0.795 0.535 0.825 0.535 0.825 0.525 1.475 0.525 1.475 0.32 1.535 0.32 1.535 0.525 1.92 0.525 1.92 0.32 1.98 0.32 1.98 0.525 2.065 0.525 ;
      POLYGON 1.915 0.705 1.875 0.705 1.875 0.75 1.86 0.75 1.86 1.18 1.8 1.18 1.8 0.705 1.795 0.705 1.795 0.645 1.915 0.645 ;
      POLYGON 1.805 2.57 1.765 2.57 1.765 3.115 1.705 3.115 1.705 2.17 1.765 2.17 1.765 2.45 1.805 2.45 ;
      POLYGON 1.775 0.465 1.715 0.465 1.715 0.255 1.33 0.255 1.33 0.465 1.27 0.465 1.27 0.195 1.775 0.195 ;
      POLYGON 1.715 0.705 1.685 0.705 1.685 1.185 1.525 1.185 1.525 1.2 1.405 1.2 1.405 1.14 1.435 1.14 1.435 1.125 1.625 1.125 1.625 0.705 1.595 0.705 1.595 0.645 1.715 0.645 ;
      POLYGON 1.32 3.115 1.26 3.115 1.26 2.6 0.98 2.6 0.98 2.54 1.26 2.54 1.26 2.185 1.32 2.185 ;
      POLYGON 0.91 3.115 0.85 3.115 0.85 2.82 0.79 2.82 0.79 2.7 0.85 2.7 0.85 1.86 0.91 1.86 ;
      POLYGON 0.64 1.525 0.37 1.525 0.37 1.465 0.58 1.465 0.58 0.32 0.64 0.32 ;
      POLYGON 0.64 2.075 0.57 2.075 0.57 3.115 0.51 3.115 0.51 2.015 0.64 2.015 ;
      RECT 0.28 0.135 0.34 1.305 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RDFFNSRQX1

MACRO RDFFNSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RDFFNSRX1 0 0 ;
  SIZE 6.2 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 5.935 1.77 5.935 2.46 5.875 2.46 5.875 1.77 5.255 1.77 5.255 2.46 5.195 2.46 5.195 1.77 1.465 1.77 1.465 2.28 1.405 2.28 1.405 1.77 0.62 1.77 0.62 2.28 0.56 2.28 0.56 1.77 0 1.77 0 1.65 0.25 1.65 0.25 1.05 0.31 1.05 0.31 1.65 1.095 1.65 1.095 1.27 1.155 1.27 1.155 1.65 1.25 1.65 1.25 1.27 1.31 1.27 1.31 1.65 1.885 1.65 1.885 1.27 1.945 1.27 1.945 1.65 5.435 1.65 5.435 1.13 5.495 1.13 5.495 1.65 5.95 1.65 5.95 1.13 6.01 1.13 6.01 1.65 6.2 1.65 ;
    END
  END VDD
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.116 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 3.580247 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 36.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 0.92 1.31 0.92 1.31 1.14 1.34 1.14 1.34 1.2 1.22 1.2 1.22 1.14 1.25 1.14 1.25 0.92 1.235 0.92 1.235 0.72 1.365 0.72 ;
    END
  END SN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 3.42 2 3.9 2.61 ;
    END
  END ExtVDD
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.27777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.415 2.69 1.565 2.825 ;
    END
  END CKN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.25 0.79 0.39 0.94 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.69295 LAYER Metal1 ;
    ANTENNADIFFAREA 3.76965 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2853 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.95425875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 152.76551 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.765 2.82 5.73 2.82 5.73 3.135 5.67 3.135 5.67 2.82 5.635 2.82 5.635 2.5 5.67 2.5 5.67 2.07 5.73 2.07 5.73 2.5 5.765 2.5 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.69295 LAYER Metal1 ;
    ANTENNADIFFAREA 3.76965 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2853 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.95425875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 152.76551 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.05 3.135 4.99 3.135 4.99 2.82 4.835 2.82 4.835 2.5 4.99 2.5 4.99 2.07 5.05 2.07 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 2.505 0.67 2.635 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 3.48 0 3.48 0 3.36 0.56 3.36 0.56 2.97 0.62 2.97 0.62 3.36 1.405 3.36 1.405 2.97 1.465 2.97 1.465 3.36 3.42 3.36 3.42 3.025 3.48 3.025 3.48 3.36 3.84 3.36 3.84 3.025 3.9 3.025 3.9 3.36 5.195 3.36 5.195 2.875 5.255 2.875 5.255 3.36 5.875 3.36 5.875 2.875 5.935 2.875 5.935 3.36 6.2 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 6.07 0.06 6.07 0.465 6.01 0.465 6.01 0.06 3.955 0.06 3.955 0.34 3.895 0.34 3.895 0.06 1.155 0.06 1.155 0.32 1.33 0.32 1.33 0.465 1.095 0.465 1.095 0.06 0.31 0.06 0.31 0.465 0.25 0.465 0.25 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.535 1.17 4.765 1.3 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.865 0.465 5.805 0.465 5.805 0.26 5.455 0.26 5.455 0.465 5.395 0.465 5.395 0.2 5.865 0.2 ;
      POLYGON 5.805 1.345 5.745 1.345 5.745 1.015 5.255 1.015 5.255 1.345 5.195 1.345 5.195 0.955 5.805 0.955 ;
      POLYGON 5.66 0.67 5.195 0.67 5.195 0.32 5.255 0.32 5.255 0.61 5.6 0.61 5.6 0.32 5.66 0.32 ;
      POLYGON 5.49 3.075 5.43 3.075 5.43 2.685 5.135 2.685 5.135 2.625 5.43 2.625 5.43 2.155 5.49 2.155 ;
      POLYGON 5.05 1.345 4.99 1.345 4.99 0.425 4.775 0.425 4.775 0.365 4.99 0.365 4.99 0.32 5.05 0.32 ;
      POLYGON 5.025 1.55 2.61 1.55 2.61 1.025 2.67 1.025 2.67 1.49 5.025 1.49 ;
      POLYGON 4.915 0.665 4.885 0.665 4.885 1.425 2.78 1.425 2.78 1.365 4.825 1.365 4.825 0.665 4.785 0.665 4.785 0.605 4.825 0.605 4.825 0.555 4.885 0.555 4.885 0.605 4.915 0.605 ;
      RECT 4.3 2.385 4.745 2.445 ;
      POLYGON 4.715 1 4.47 1 4.47 0.25 4.46 0.25 4.46 0.23 4.445 0.23 4.445 0.17 4.46 0.17 4.46 0.13 4.52 0.13 4.52 0.17 4.53 0.17 4.53 0.94 4.715 0.94 ;
      RECT 4.65 0.135 4.71 0.84 ;
      POLYGON 4.39 1.22 4.38 1.22 4.38 1.25 4.32 1.25 4.32 1.22 4.2 1.22 4.2 1.255 4.14 1.255 4.14 1.13 4.2 1.13 4.2 1.16 4.32 1.16 4.32 1.13 4.33 1.13 4.33 0.415 4.2 0.415 4.2 0.47 3.715 0.47 3.715 0.3 3.6 0.3 3.6 0.24 3.775 0.24 3.775 0.41 4.14 0.41 4.14 0.32 4.2 0.32 4.2 0.355 4.39 0.355 ;
      POLYGON 4.245 0.65 4.185 0.65 4.185 0.615 3.735 0.615 3.735 0.65 3.615 0.65 3.615 0.59 3.675 0.59 3.675 0.555 4.185 0.555 4.185 0.53 4.245 0.53 ;
      POLYGON 4.245 0.89 4.185 0.89 4.185 0.86 3.85 0.86 3.85 0.8 4.185 0.8 4.185 0.77 4.245 0.77 ;
      POLYGON 4.21 3.17 4.15 3.17 4.15 2.78 3.35 2.78 3.35 2.72 4.15 2.72 4.15 2 4.21 2 ;
      POLYGON 4.005 2.93 3.275 2.93 3.275 3.17 3.215 3.17 3.215 2 3.275 2 3.275 2.87 4.005 2.87 ;
      RECT 3.74 1.13 3.995 1.25 ;
      POLYGON 3.655 1.25 3.42 1.25 3.42 0.32 3.48 0.32 3.48 1.19 3.595 1.19 3.595 1.13 3.655 1.13 ;
      POLYGON 3.275 1.255 3.215 1.255 3.215 0.65 2.39 0.65 2.39 1.485 2.33 1.485 2.33 0.32 2.39 0.32 2.39 0.59 3.155 0.59 3.155 0.58 3.215 0.58 3.215 0.32 3.275 0.32 ;
      POLYGON 2.27 1.19 2.185 1.19 2.185 1.485 2.125 1.485 2.125 1.13 2.21 1.13 2.21 0.585 1.515 0.585 1.515 1.27 1.635 1.27 1.635 1.485 1.455 1.485 1.455 0.585 1.12 0.585 1.12 0.595 1.09 0.595 1.09 1.14 1.12 1.14 1.12 1.2 1 1.2 1 1.14 1.03 1.14 1.03 0.595 1 0.595 1 0.535 1.03 0.535 1.03 0.525 1.68 0.525 1.68 0.32 1.74 0.32 1.74 0.525 2.125 0.525 2.125 0.32 2.185 0.32 2.185 0.525 2.27 0.525 ;
      POLYGON 2.12 0.705 2.08 0.705 2.08 0.75 2.065 0.75 2.065 1.18 2.005 1.18 2.005 0.705 2 0.705 2 0.645 2.12 0.645 ;
      POLYGON 1.98 0.465 1.92 0.465 1.92 0.255 1.535 0.255 1.535 0.465 1.475 0.465 1.475 0.195 1.98 0.195 ;
      POLYGON 1.92 0.705 1.89 0.705 1.89 1.185 1.61 1.185 1.61 1.125 1.83 1.125 1.83 0.705 1.8 0.705 1.8 0.645 1.92 0.645 ;
      POLYGON 1.73 3.03 1.67 3.03 1.67 3.115 1.61 3.115 1.61 2.97 1.67 2.97 1.67 2.605 1.3 2.605 1.3 2.545 1.67 2.545 1.67 2.28 1.61 2.28 1.61 2.065 1.67 2.065 1.67 2.13 1.73 2.13 ;
      POLYGON 1.26 2.39 1.15 2.39 1.15 2.97 1.26 2.97 1.26 3.115 1.2 3.115 1.2 3.03 1.09 3.03 1.09 2.33 1.2 2.33 1.2 1.985 1.125 1.985 1.125 1.925 1.26 1.925 ;
      POLYGON 0.93 3.115 0.87 3.115 0.87 2.435 0.345 2.435 0.345 2.375 0.87 2.375 0.87 2.065 0.93 2.065 ;
      POLYGON 0.845 1.485 0.435 1.485 0.435 1.56 0.375 1.56 0.375 1.425 0.785 1.425 0.785 0.32 0.845 0.32 ;
      RECT 0.615 0.135 0.675 1.305 ;
      POLYGON 0.555 0.985 0.515 0.985 0.515 1.265 0.455 1.265 0.455 0.32 0.515 0.32 0.515 0.865 0.555 0.865 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RDFFNSRX1

MACRO RDFFNSX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RDFFNSX1 0 0 ;
  SIZE 5.8 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 1.77 5.53 1.77 5.53 2.46 5.47 2.46 5.47 1.77 4.85 1.77 4.85 2.46 4.79 2.46 4.79 1.77 1.115 1.77 1.115 2.4 1.055 2.4 1.055 1.77 0.26 1.77 0.26 2.4 0.2 2.4 0.2 1.77 -0.005 1.77 -0.005 1.65 0.7 1.65 0.7 1.165 0.76 1.165 0.76 1.65 1.38 1.65 1.38 1.25 1.385 1.25 1.385 1.165 1.445 1.165 1.445 1.38 1.44 1.38 1.44 1.65 5.03 1.65 5.03 1.13 5.09 1.13 5.09 1.65 5.44 1.65 5.44 1.13 5.5 1.13 5.5 1.65 5.8 1.65 ;
    END
  END VDD
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0516 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.5925925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 21.9444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.965 1.095 0.81 1.095 0.81 1.035 0.84 1.035 0.84 0.72 0.9 0.72 0.9 0.79 0.965 0.79 ;
    END
  END SN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.495 2.61 3.015 2.61 3.015 2 3.145 2 3.145 1.89 3.395 1.89 3.395 2 3.495 2 ;
    END
  END ExtVDD
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.64814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 2.69 1.185 2.845 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.86725 LAYER Metal1 ;
    ANTENNADIFFAREA 3.6343 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2529 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.24574925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 138.76631075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.365 2.82 5.325 2.82 5.325 3.135 5.265 3.135 5.265 2.82 5.235 2.82 5.235 2.5 5.265 2.5 5.265 2.07 5.325 2.07 5.325 2.5 5.365 2.5 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.86725 LAYER Metal1 ;
    ANTENNADIFFAREA 3.6343 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2529 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.24574925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 138.76631075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.645 3.135 4.585 3.135 4.585 2.82 4.435 2.82 4.435 2.5 4.585 2.5 4.585 2.07 4.645 2.07 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.462963 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.2 2.5 0.365 2.63 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 3.48 0 3.48 0 3.36 0.2 3.36 0.2 2.97 0.26 2.97 0.26 3.36 1.055 3.36 1.055 2.97 1.115 2.97 1.115 3.36 3.015 3.36 3.015 3.025 3.075 3.025 3.075 3.36 3.435 3.36 3.435 3.025 3.495 3.025 3.495 3.36 4.79 3.36 4.79 2.875 4.85 2.875 4.85 3.36 5.47 3.36 5.47 2.875 5.53 2.875 5.53 3.36 5.8 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 0.06 5.5 0.06 5.5 0.465 5.44 0.465 5.44 0.06 3.59 0.06 3.59 0.465 3.53 0.465 3.53 0.06 0.76 0.06 0.76 0.32 0.935 0.32 0.935 0.465 0.7 0.465 0.7 0.06 0 0.06 0 -0.06 5.8 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.537037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.365 1.525 4.055 1.525 4.055 1.37 3.91 1.37 3.91 0.41 3.97 0.41 3.97 1.31 4.365 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.295 1.345 5.235 1.345 5.235 1.015 4.85 1.015 4.85 1.345 4.79 1.345 4.79 0.955 5.295 0.955 ;
      POLYGON 5.19 0.465 5.13 0.465 5.13 0.42 4.85 0.42 4.85 0.495 4.79 0.495 4.79 0.32 4.85 0.32 4.85 0.36 5.13 0.36 5.13 0.32 5.19 0.32 ;
      POLYGON 5.085 3.08 5.025 3.08 5.025 2.655 4.73 2.655 4.73 2.595 5.025 2.595 5.025 2.16 5.085 2.16 ;
      RECT 4.585 0.32 4.645 1.345 ;
      RECT 3.895 2.385 4.34 2.445 ;
      POLYGON 4.335 1.13 4.065 1.13 4.065 0.25 4.055 0.25 4.055 0.23 4.04 0.23 4.04 0.17 4.055 0.17 4.055 0.13 4.115 0.13 4.115 0.17 4.125 0.17 4.125 1.07 4.335 1.07 ;
      RECT 4.245 0.135 4.305 0.995 ;
      POLYGON 3.995 1.51 3.735 1.51 3.735 0.83 3.2 0.83 3.2 0.245 3.26 0.245 3.26 0.77 3.735 0.77 3.735 0.32 3.795 0.32 3.795 1.45 3.995 1.45 ;
      POLYGON 3.805 3.17 3.745 3.17 3.745 2.78 2.945 2.78 2.945 2.72 3.745 2.72 3.745 2 3.805 2 ;
      POLYGON 3.6 2.93 2.87 2.93 2.87 3.17 2.81 3.17 2.81 2 2.87 2 2.87 2.87 3.6 2.87 ;
      RECT 3.31 1.24 3.59 1.525 ;
      RECT 3.015 0.32 3.075 1.455 ;
      POLYGON 2.87 1.52 2.58 1.52 2.58 1.46 2.81 1.46 2.81 0.32 2.87 0.32 ;
      RECT 2.275 0.6 2.335 1.18 ;
      POLYGON 1.95 0.83 1.89 0.83 1.89 1.38 1.83 1.38 1.83 0.32 1.89 0.32 1.89 0.77 1.95 0.77 ;
      POLYGON 1.685 1.38 1.625 1.38 1.625 0.585 1.12 0.585 1.12 1.165 1.24 1.165 1.24 1.38 0.905 1.38 0.905 1.165 1.06 1.165 1.06 0.585 0.725 0.585 0.725 0.595 0.695 0.595 0.695 1.035 0.725 1.035 0.725 1.095 0.605 1.095 0.605 1.035 0.635 1.035 0.635 0.595 0.605 0.595 0.605 0.535 0.635 0.535 0.635 0.525 1.185 0.525 1.185 0.32 1.245 0.32 1.245 0.525 1.625 0.525 1.625 0.32 1.685 0.32 ;
      POLYGON 1.335 0.705 1.305 0.705 1.305 1.035 1.335 1.035 1.335 1.095 1.215 1.095 1.215 1.035 1.245 1.035 1.245 0.705 1.215 0.705 1.215 0.645 1.335 0.645 ;
      POLYGON 1.32 3.115 1.26 3.115 1.26 2.6 0.98 2.6 0.98 2.54 1.26 2.54 1.26 2.185 1.32 2.185 ;
      POLYGON 0.91 3.115 0.85 3.115 0.85 2.82 0.79 2.82 0.79 2.7 0.85 2.7 0.85 1.86 0.91 1.86 ;
      POLYGON 0.64 2.1 0.57 2.1 0.57 3.115 0.51 3.115 0.51 2.015 0.61 2.015 0.61 2.04 0.64 2.04 ;
      POLYGON 0.45 1.52 0.29 1.52 0.29 1.46 0.39 1.46 0.39 0.32 0.45 0.32 ;
      RECT 0.1 0.135 0.16 1.2 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RDFFNSX1

MACRO RDFFNX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RDFFNX1 0 0 ;
  SIZE 5.2 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.2 1.77 4.93 1.77 4.93 2.46 4.87 2.46 4.87 1.77 4.255 1.77 4.255 2.465 4.195 2.465 4.195 1.77 1.035 1.77 1.035 2.4 0.975 2.4 0.975 1.77 0.255 1.77 0.255 2.4 0.195 2.4 0.195 1.77 0 1.77 0 1.65 0.895 1.65 0.895 1.11 0.955 1.11 0.955 1.65 4.3 1.65 4.3 1.13 4.36 1.13 4.36 1.65 5.2 1.65 ;
    END
  END VDD
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.29615 LAYER Metal1 ;
    ANTENNADIFFAREA 3.206275 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2529 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.9875445 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 122.08778175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.05 3.13 3.99 3.13 3.99 2.82 3.835 2.82 3.835 2.5 3.99 2.5 3.99 2.075 4.05 2.075 ;
    END
  END QN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.9 2.61 2.42 2.61 2.42 2 2.57 2 2.57 1.89 2.82 1.89 2.82 2 2.9 2 ;
    END
  END ExtVDD
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.29615 LAYER Metal1 ;
    ANTENNADIFFAREA 3.206275 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2529 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.9875445 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 122.08778175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.765 2.82 4.725 2.82 4.725 3.135 4.665 3.135 4.665 2.82 4.635 2.82 4.635 2.5 4.665 2.5 4.665 2.07 4.725 2.07 4.725 2.5 4.765 2.5 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.185 2.69 0.365 2.83 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.2 3.48 0 3.48 0 3.36 0.195 3.36 0.195 2.97 0.255 2.97 0.255 3.36 0.975 3.36 0.975 2.97 1.035 2.97 1.035 3.36 2.42 3.36 2.42 3.025 2.48 3.025 2.48 3.36 2.84 3.36 2.84 3.025 2.9 3.025 2.9 3.36 4.195 3.36 4.195 2.87 4.255 2.87 4.255 3.36 4.87 3.36 4.87 2.875 4.93 2.875 4.93 3.36 5.2 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.2 0.06 4.36 0.06 4.36 0.465 4.3 0.465 4.3 0.06 2.995 0.06 2.995 0.625 2.935 0.625 2.935 0.06 0.955 0.06 0.955 0.54 0.895 0.54 0.895 0.06 0 0.06 0 -0.06 5.2 -0.06 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.985 2.475 1.165 2.63 ;
    END
  END CKN
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0441 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.361111 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 17.68518525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.435 1.17 3.565 1.36 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 4.49 3.075 4.43 3.075 4.43 2.685 4.135 2.685 4.135 2.625 4.43 2.625 4.43 2.165 4.49 2.165 ;
      POLYGON 4.05 1.345 3.99 1.345 3.99 1.05 3.96 1.05 3.96 0.93 3.99 0.93 3.99 0.32 4.05 0.32 ;
      RECT 3.775 0.14 3.835 1.45 ;
      RECT 3.3 2.615 3.745 2.675 ;
      POLYGON 3.42 1.525 3.14 1.525 3.14 1.025 2.66 1.025 2.66 0.38 2.72 0.38 2.72 0.965 3.14 0.965 3.14 0.48 3.2 0.48 3.2 1.465 3.42 1.465 ;
      RECT 3.31 0.48 3.37 1.215 ;
      POLYGON 3.21 3.17 3.15 3.17 3.15 2.78 2.35 2.78 2.35 2.72 3.15 2.72 3.15 2 3.21 2 ;
      POLYGON 3.005 2.93 2.275 2.93 2.275 3.17 2.215 3.17 2.215 2 2.275 2 2.275 2.87 3.005 2.87 ;
      POLYGON 2.995 1.555 2.735 1.555 2.735 1.26 2.935 1.26 2.935 1.255 2.995 1.255 ;
      RECT 2.42 0.48 2.48 1.47 ;
      POLYGON 2.275 1.54 2.005 1.54 2.005 1.48 2.215 1.48 2.215 0.48 2.275 0.48 ;
      POLYGON 2.125 1.02 2.005 1.02 2.005 0.96 2.035 0.96 2.035 0.86 1.365 0.86 1.365 1.325 1.305 1.325 1.305 0.38 1.365 0.38 1.365 0.8 2.095 0.8 2.095 0.96 2.125 0.96 ;
      POLYGON 1.3 3.03 1.24 3.03 1.24 3.115 1.18 3.115 1.18 2.97 1.24 2.97 1.24 2.795 0.895 2.795 0.895 2.735 1.24 2.735 1.24 2.4 1.18 2.4 1.18 2.185 1.24 2.185 1.24 2.25 1.3 2.25 ;
      POLYGON 1.16 1.325 1.1 1.325 1.1 0.85 0.89 0.85 0.89 0.98 0.92 0.98 0.92 1.04 0.8 1.04 0.8 0.98 0.83 0.98 0.83 0.67 0.8 0.67 0.8 0.61 0.92 0.61 0.92 0.67 0.89 0.67 0.89 0.79 1.1 0.79 1.1 0.395 1.16 0.395 ;
      POLYGON 0.83 3.115 0.77 3.115 0.77 2.795 0.68 2.795 0.68 2.735 0.77 2.735 0.77 1.885 0.83 1.885 ;
      POLYGON 0.645 1.325 0.635 1.325 0.635 1.525 0.475 1.525 0.475 1.465 0.575 1.465 0.575 1.11 0.585 1.11 0.585 0.395 0.645 0.395 ;
      POLYGON 0.61 2.155 0.565 2.155 0.565 3.115 0.505 3.115 0.505 2.095 0.55 2.095 0.55 1.84 0.61 1.84 ;
      RECT 0.305 0.145 0.365 1.545 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RDFFNX1

MACRO RDFFQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RDFFQX1 0 0 ;
  SIZE 4.6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.77 4.37 1.77 4.37 2.465 4.31 2.465 4.31 1.77 1.04 1.77 1.04 2.405 0.98 2.405 0.98 1.77 0.26 1.77 0.26 2.405 0.2 2.405 0.2 1.77 0 1.77 0 1.65 0.9 1.65 0.9 1.115 0.96 1.115 0.96 1.65 4.305 1.65 4.305 1.135 4.365 1.135 4.365 1.65 4.6 1.65 ;
    END
  END VDD
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.388889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.965 2.505 1.165 2.65 ;
    END
  END CK
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.905 2.615 2.425 2.615 2.425 2.005 2.575 2.005 2.575 1.895 2.825 1.895 2.825 2.005 2.905 2.005 ;
    END
  END ExtVDD
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.79195 LAYER Metal1 ;
    ANTENNADIFFAREA 2.739875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20745 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.2788625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 131.97396975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.17 2.825 4.165 2.825 4.165 3.14 4.105 3.14 4.105 2.825 4.04 2.825 4.04 2.695 4.105 2.695 4.105 2.075 4.165 2.075 4.165 2.695 4.17 2.695 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.19 2.695 0.37 2.84 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 3.48 0 3.48 0 3.36 0.2 3.36 0.2 2.975 0.26 2.975 0.26 3.36 0.98 3.36 0.98 2.975 1.04 2.975 1.04 3.36 2.425 3.36 2.425 3.03 2.485 3.03 2.485 3.36 2.845 3.36 2.845 3.03 2.905 3.03 2.905 3.36 4.31 3.36 4.31 2.88 4.37 2.88 4.37 3.36 4.6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 0.06 4.365 0.06 4.365 0.47 4.305 0.47 4.305 0.06 3 0.06 3 0.63 2.94 0.63 2.94 0.06 0.96 0.06 0.96 0.545 0.9 0.545 0.9 0.06 0 0.06 0 -0.06 4.6 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0441 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.361111 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 17.962963 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.44 1.175 3.6 1.365 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 4.055 1.35 3.995 1.35 3.995 1.055 3.965 1.055 3.965 0.935 3.995 0.935 3.995 0.325 4.055 0.325 ;
      RECT 3.78 0.145 3.84 1.455 ;
      RECT 3.305 2.62 3.75 2.68 ;
      POLYGON 3.425 1.53 3.145 1.53 3.145 1.03 2.665 1.03 2.665 0.385 2.725 0.385 2.725 0.97 3.145 0.97 3.145 0.485 3.205 0.485 3.205 1.47 3.425 1.47 ;
      RECT 3.315 0.485 3.375 1.22 ;
      POLYGON 3.215 3.175 3.155 3.175 3.155 2.785 2.355 2.785 2.355 2.725 3.155 2.725 3.155 2.005 3.215 2.005 ;
      POLYGON 3.01 2.935 2.28 2.935 2.28 3.175 2.22 3.175 2.22 2.005 2.28 2.005 2.28 2.875 3.01 2.875 ;
      POLYGON 3 1.56 2.74 1.56 2.74 1.265 2.94 1.265 2.94 1.26 3 1.26 ;
      RECT 2.425 0.485 2.485 1.475 ;
      POLYGON 2.28 1.545 2.01 1.545 2.01 1.485 2.22 1.485 2.22 0.485 2.28 0.485 ;
      POLYGON 2.13 1.025 2.01 1.025 2.01 0.965 2.04 0.965 2.04 0.865 1.37 0.865 1.37 1.33 1.31 1.33 1.31 0.385 1.37 0.385 1.37 0.805 2.1 0.805 2.1 0.965 2.13 0.965 ;
      POLYGON 1.305 3.035 1.245 3.035 1.245 3.12 1.185 3.12 1.185 2.975 1.245 2.975 1.245 2.8 0.9 2.8 0.9 2.74 1.245 2.74 1.245 2.405 1.185 2.405 1.185 2.19 1.245 2.19 1.245 2.255 1.305 2.255 ;
      POLYGON 1.165 1.33 1.105 1.33 1.105 0.855 0.895 0.855 0.895 0.985 0.925 0.985 0.925 1.045 0.805 1.045 0.805 0.985 0.835 0.985 0.835 0.675 0.805 0.675 0.805 0.615 0.925 0.615 0.925 0.675 0.895 0.675 0.895 0.795 1.105 0.795 1.105 0.4 1.165 0.4 ;
      POLYGON 0.835 3.12 0.775 3.12 0.775 2.61 0.69 2.61 0.69 2.55 0.775 2.55 0.775 2.19 0.835 2.19 ;
      POLYGON 0.65 1.33 0.64 1.33 0.64 1.53 0.48 1.53 0.48 1.47 0.58 1.47 0.58 1.115 0.59 1.115 0.59 0.4 0.65 0.4 ;
      POLYGON 0.615 2.16 0.57 2.16 0.57 3.12 0.51 3.12 0.51 2.1 0.555 2.1 0.555 1.845 0.615 1.845 ;
      RECT 0.31 0.15 0.37 1.55 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RDFFQX1

MACRO RDFFRQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RDFFRQX1 0 0 ;
  SIZE 5.6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 5.185 1.77 5.185 2.46 5.125 2.46 5.125 1.77 1.56 1.77 1.56 2.385 1.5 2.385 1.5 1.77 1.115 1.77 1.115 2.4 1.055 2.4 1.055 1.77 0.26 1.77 0.26 2.4 0.2 2.4 0.2 1.77 -0.005 1.77 -0.005 1.65 0.89 1.65 0.89 1.27 0.95 1.27 0.95 1.65 1.44 1.65 1.44 1.27 1.5 1.27 1.5 1.65 5.03 1.65 5.03 1.13 5.09 1.13 5.09 1.65 5.6 1.65 ;
    END
  END VDD
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.495 2.61 3.015 2.61 3.015 2 3.145 2 3.145 1.89 3.395 1.89 3.395 2 3.495 2 ;
    END
  END ExtVDD
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.64 2.59 1.63 2.59 1.63 2.63 1.435 2.63 1.435 2.5 1.63 2.5 1.63 2.53 1.64 2.53 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5387 LAYER Metal1 ;
    ANTENNADIFFAREA 3.382925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.23985 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.923077 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 137.64853025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.98 3.135 4.92 3.135 4.92 2.82 4.835 2.82 4.835 2.5 4.92 2.5 4.92 2.07 4.98 2.07 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.5555555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.195 2.5 0.365 2.63 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 3.48 0 3.48 0 3.36 0.2 3.36 0.2 2.97 0.26 2.97 0.26 3.36 1.055 3.36 1.055 2.97 1.115 2.97 1.115 3.36 1.5 3.36 1.5 2.97 1.56 2.97 1.56 3.36 3.015 3.36 3.015 3.025 3.075 3.025 3.075 3.36 3.435 3.36 3.435 3.025 3.495 3.025 3.495 3.36 5.125 3.36 5.125 2.875 5.185 2.875 5.185 3.36 5.6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5.46 0.06 5.46 0.465 5.4 0.465 5.4 0.06 5.05 0.06 5.05 0.465 4.99 0.465 4.99 0.06 3.59 0.06 3.59 0.465 3.53 0.465 3.53 0.06 1.405 0.06 1.405 0.465 1.345 0.465 1.345 0.06 0.95 0.06 0.95 0.465 0.89 0.465 0.89 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.83333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.025 2.69 1.185 2.845 ;
    END
  END CK
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.537037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.365 1.525 4.055 1.525 4.055 1.37 3.91 1.37 3.91 0.41 3.97 0.41 3.97 1.31 4.365 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.4 1.345 5.34 1.345 5.34 1.015 4.85 1.015 4.85 1.345 4.79 1.345 4.79 0.955 5.4 0.955 ;
      POLYGON 5.255 0.67 4.79 0.67 4.79 0.32 4.85 0.32 4.85 0.61 5.195 0.61 5.195 0.32 5.255 0.32 ;
      RECT 4.585 0.32 4.645 1.345 ;
      RECT 3.895 2.385 4.34 2.445 ;
      POLYGON 4.335 1.08 4.065 1.08 4.065 0.25 4.055 0.25 4.055 0.23 4.04 0.23 4.04 0.17 4.055 0.17 4.055 0.13 4.115 0.13 4.115 0.17 4.125 0.17 4.125 1.02 4.335 1.02 ;
      POLYGON 3.995 1.51 3.735 1.51 3.735 0.685 3.2 0.685 3.2 0.52 3.26 0.52 3.26 0.625 3.735 0.625 3.735 0.32 3.795 0.32 3.795 1.45 3.995 1.45 ;
      POLYGON 3.805 3.17 3.745 3.17 3.745 2.78 2.945 2.78 2.945 2.72 3.745 2.72 3.745 2 3.805 2 ;
      POLYGON 3.6 2.93 2.87 2.93 2.87 3.17 2.81 3.17 2.81 2 2.87 2 2.87 2.87 3.6 2.87 ;
      RECT 3.31 1.24 3.59 1.525 ;
      RECT 3.015 0.32 3.075 1.455 ;
      POLYGON 2.87 1.52 2.58 1.52 2.58 1.46 2.81 1.46 2.81 0.32 2.87 0.32 ;
      RECT 2.275 0.71 2.335 1.285 ;
      POLYGON 1.945 1.485 1.885 1.485 1.885 0.85 1.755 0.85 1.755 0.32 1.815 0.32 1.815 0.79 1.945 0.79 ;
      POLYGON 1.805 2.57 1.765 2.57 1.765 3.115 1.705 3.115 1.705 2.17 1.765 2.17 1.765 2.45 1.805 2.45 ;
      POLYGON 1.74 1.485 1.68 1.485 1.68 1.2 1.19 1.2 1.19 1.485 1.13 1.485 1.13 1.2 0.795 1.2 0.795 1.14 1.28 1.14 1.28 0.595 0.795 0.595 0.795 0.535 1.095 0.535 1.095 0.32 1.155 0.32 1.155 0.535 1.55 0.535 1.55 0.32 1.61 0.32 1.61 0.595 1.34 0.595 1.34 1.14 1.74 1.14 ;
      POLYGON 1.32 3.115 1.26 3.115 1.26 2.6 0.98 2.6 0.98 2.54 1.26 2.54 1.26 2.185 1.32 2.185 ;
      POLYGON 0.91 3.115 0.85 3.115 0.85 2.64 0.79 2.64 0.79 2.52 0.85 2.52 0.85 2.185 0.91 2.185 ;
      POLYGON 0.64 1.525 0.37 1.525 0.37 1.465 0.58 1.465 0.58 0.32 0.64 0.32 ;
      POLYGON 0.64 2.075 0.57 2.075 0.57 3.115 0.51 3.115 0.51 2.015 0.64 2.015 ;
      RECT 0.28 0.135 0.34 1.305 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RDFFRQX1

MACRO RDFFRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RDFFRX1 0 0 ;
  SIZE 5.8 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 1.77 5.53 1.77 5.53 2.46 5.47 2.46 5.47 1.77 4.85 1.77 4.85 2.46 4.79 2.46 4.79 1.77 1.56 1.77 1.56 2.385 1.5 2.385 1.5 1.77 1.115 1.77 1.115 2.4 1.055 2.4 1.055 1.77 0.26 1.77 0.26 2.4 0.2 2.4 0.2 1.77 -0.005 1.77 -0.005 1.65 0.89 1.65 0.89 1.27 0.95 1.27 0.95 1.65 1.44 1.65 1.44 1.27 1.5 1.27 1.5 1.65 5.03 1.65 5.03 1.13 5.09 1.13 5.09 1.65 5.8 1.65 ;
    END
  END VDD
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.495 2.61 3.015 2.61 3.015 2 3.145 2 3.145 1.89 3.395 1.89 3.395 2 3.495 2 ;
    END
  END ExtVDD
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.4074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.64 2.59 1.63 2.59 1.63 2.65 1.435 2.65 1.435 2.455 1.63 2.455 1.63 2.53 1.64 2.53 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.86085 LAYER Metal1 ;
    ANTENNADIFFAREA 3.681325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2853 LAYER Metal1 ;
      ANTENNAMAXAREACAR 17.03767975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 124.7844375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.365 2.82 5.325 2.82 5.325 3.135 5.265 3.135 5.265 2.82 5.235 2.82 5.235 2.505 5.265 2.505 5.265 2.07 5.325 2.07 5.325 2.505 5.365 2.505 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.86085 LAYER Metal1 ;
    ANTENNADIFFAREA 3.681325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2853 LAYER Metal1 ;
      ANTENNAMAXAREACAR 17.03767975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 124.7844375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.645 3.135 4.585 3.135 4.585 2.82 4.435 2.82 4.435 2.5 4.585 2.5 4.585 2.07 4.645 2.07 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.16 2.5 0.365 2.63 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 3.48 0 3.48 0 3.36 0.2 3.36 0.2 2.97 0.26 2.97 0.26 3.36 1.055 3.36 1.055 2.97 1.115 2.97 1.115 3.36 1.5 3.36 1.5 2.97 1.56 2.97 1.56 3.36 3.015 3.36 3.015 3.025 3.075 3.025 3.075 3.36 3.435 3.36 3.435 3.025 3.495 3.025 3.495 3.36 4.79 3.36 4.79 2.875 4.85 2.875 4.85 3.36 5.47 3.36 5.47 2.875 5.53 2.875 5.53 3.36 5.8 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 0.06 5.46 0.06 5.46 0.465 5.4 0.465 5.4 0.06 5.05 0.06 5.05 0.465 4.99 0.465 4.99 0.06 3.59 0.06 3.59 0.465 3.53 0.465 3.53 0.06 1.405 0.06 1.405 0.465 1.345 0.465 1.345 0.06 0.95 0.06 0.95 0.465 0.89 0.465 0.89 0.06 0 0.06 0 -0.06 5.8 -0.06 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.83333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.025 2.69 1.185 2.845 ;
    END
  END CK
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.62962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.375 1.525 4.055 1.525 4.055 1.37 3.91 1.37 3.91 0.41 3.97 0.41 3.97 1.31 4.375 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.4 1.345 5.34 1.345 5.34 1.015 4.85 1.015 4.85 1.345 4.79 1.345 4.79 0.955 5.4 0.955 ;
      POLYGON 5.255 0.67 4.79 0.67 4.79 0.32 4.85 0.32 4.85 0.61 5.195 0.61 5.195 0.32 5.255 0.32 ;
      POLYGON 5.085 3.075 5.025 3.075 5.025 2.68 4.73 2.68 4.73 2.62 5.025 2.62 5.025 2.155 5.085 2.155 ;
      RECT 4.585 0.32 4.645 1.345 ;
      RECT 3.895 2.385 4.34 2.445 ;
      POLYGON 4.335 1.08 4.065 1.08 4.065 0.25 4.055 0.25 4.055 0.23 4.04 0.23 4.04 0.17 4.055 0.17 4.055 0.13 4.115 0.13 4.115 0.17 4.125 0.17 4.125 1.02 4.335 1.02 ;
      POLYGON 3.995 1.51 3.735 1.51 3.735 0.685 3.2 0.685 3.2 0.52 3.26 0.52 3.26 0.625 3.735 0.625 3.735 0.32 3.795 0.32 3.795 1.45 3.995 1.45 ;
      POLYGON 3.805 3.17 3.745 3.17 3.745 2.78 2.945 2.78 2.945 2.72 3.745 2.72 3.745 2 3.805 2 ;
      POLYGON 3.6 2.93 2.87 2.93 2.87 3.17 2.81 3.17 2.81 2 2.87 2 2.87 2.87 3.6 2.87 ;
      RECT 3.31 1.24 3.59 1.525 ;
      RECT 3.015 0.32 3.075 1.455 ;
      POLYGON 2.87 1.52 2.58 1.52 2.58 1.46 2.81 1.46 2.81 0.32 2.87 0.32 ;
      RECT 2.275 0.71 2.335 1.285 ;
      POLYGON 1.945 1.485 1.885 1.485 1.885 0.85 1.755 0.85 1.755 0.32 1.815 0.32 1.815 0.79 1.945 0.79 ;
      POLYGON 1.805 2.57 1.765 2.57 1.765 3.115 1.705 3.115 1.705 2.17 1.765 2.17 1.765 2.45 1.805 2.45 ;
      POLYGON 1.74 1.485 1.68 1.485 1.68 1.2 1.19 1.2 1.19 1.485 1.13 1.485 1.13 1.2 0.795 1.2 0.795 1.14 1.28 1.14 1.28 0.595 0.795 0.595 0.795 0.535 1.095 0.535 1.095 0.32 1.155 0.32 1.155 0.535 1.55 0.535 1.55 0.32 1.61 0.32 1.61 0.595 1.34 0.595 1.34 1.14 1.74 1.14 ;
      POLYGON 1.32 3.115 1.26 3.115 1.26 2.6 0.98 2.6 0.98 2.54 1.26 2.54 1.26 2.185 1.32 2.185 ;
      POLYGON 0.91 3.115 0.85 3.115 0.85 2.625 0.79 2.625 0.79 2.505 0.85 2.505 0.85 2.185 0.91 2.185 ;
      POLYGON 0.64 1.525 0.37 1.525 0.37 1.465 0.58 1.465 0.58 0.32 0.64 0.32 ;
      POLYGON 0.64 2.075 0.57 2.075 0.57 3.115 0.51 3.115 0.51 2.015 0.64 2.015 ;
      RECT 0.28 0.135 0.34 1.305 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RDFFRX1

MACRO RDFFSQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RDFFSQX1 0 0 ;
  SIZE 5.6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 5.425 1.77 5.425 2.46 5.365 2.46 5.365 1.77 1.115 1.77 1.115 2.4 1.055 2.4 1.055 1.77 0.26 1.77 0.26 2.4 0.2 2.4 0.2 1.77 -0.005 1.77 -0.005 1.65 0.7 1.65 0.7 1.165 0.76 1.165 0.76 1.65 1.38 1.65 1.38 1.25 1.385 1.25 1.385 1.165 1.445 1.165 1.445 1.38 1.44 1.38 1.44 1.65 5.03 1.65 5.03 1.13 5.09 1.13 5.09 1.65 5.44 1.65 5.44 1.13 5.5 1.13 5.5 1.65 5.6 1.65 ;
    END
  END VDD
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.08745 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.699074 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 27.5925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.37 0.54 4.305 0.54 4.305 0.995 4.245 0.995 4.245 0.54 4.235 0.54 4.235 0.41 4.245 0.41 4.245 0.135 4.305 0.135 4.305 0.41 4.37 0.41 ;
    END
  END SN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.495 2.61 3.015 2.61 3.015 2 3.145 2 3.145 1.89 3.395 1.89 3.395 2 3.495 2 ;
    END
  END ExtVDD
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.53805 LAYER Metal1 ;
    ANTENNADIFFAREA 3.3359 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20745 LAYER Metal1 ;
      ANTENNAMAXAREACAR 21.87539175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 155.878525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.22 3.135 5.16 3.135 5.16 2.82 5.035 2.82 5.035 2.5 5.16 2.5 5.16 2.07 5.22 2.07 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.015 2.69 1.185 2.845 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.16 2.5 0.365 2.63 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 3.48 0 3.48 0 3.36 0.2 3.36 0.2 2.97 0.26 2.97 0.26 3.36 1.055 3.36 1.055 2.97 1.115 2.97 1.115 3.36 3.015 3.36 3.015 3.025 3.075 3.025 3.075 3.36 3.435 3.36 3.435 3.025 3.495 3.025 3.495 3.36 5.365 3.36 5.365 2.875 5.425 2.875 5.425 3.36 5.6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5.5 0.06 5.5 0.465 5.44 0.465 5.44 0.06 3.59 0.06 3.59 0.465 3.53 0.465 3.53 0.06 0.76 0.06 0.76 0.32 0.935 0.32 0.935 0.465 0.7 0.465 0.7 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.537037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.365 1.525 4.055 1.525 4.055 1.37 3.91 1.37 3.91 0.41 3.97 0.41 3.97 1.31 4.365 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.295 1.345 5.235 1.345 5.235 1.015 4.85 1.015 4.85 1.345 4.79 1.345 4.79 0.955 5.295 0.955 ;
      POLYGON 5.19 0.465 5.13 0.465 5.13 0.42 4.85 0.42 4.85 0.495 4.79 0.495 4.79 0.32 4.85 0.32 4.85 0.36 5.13 0.36 5.13 0.32 5.19 0.32 ;
      RECT 4.585 0.32 4.645 1.345 ;
      RECT 3.895 2.385 4.34 2.445 ;
      POLYGON 4.335 1.13 4.065 1.13 4.065 0.25 4.055 0.25 4.055 0.23 4.04 0.23 4.04 0.17 4.055 0.17 4.055 0.13 4.115 0.13 4.115 0.17 4.125 0.17 4.125 1.07 4.335 1.07 ;
      POLYGON 3.995 1.51 3.735 1.51 3.735 0.83 3.2 0.83 3.2 0.245 3.26 0.245 3.26 0.77 3.735 0.77 3.735 0.32 3.795 0.32 3.795 1.45 3.995 1.45 ;
      POLYGON 3.805 3.17 3.745 3.17 3.745 2.78 2.945 2.78 2.945 2.72 3.745 2.72 3.745 2 3.805 2 ;
      POLYGON 3.6 2.93 2.87 2.93 2.87 3.17 2.81 3.17 2.81 2 2.87 2 2.87 2.87 3.6 2.87 ;
      RECT 3.31 1.24 3.59 1.525 ;
      RECT 3.015 0.32 3.075 1.455 ;
      POLYGON 2.87 1.52 2.58 1.52 2.58 1.46 2.81 1.46 2.81 0.32 2.87 0.32 ;
      RECT 2.275 0.6 2.335 1.18 ;
      POLYGON 1.95 0.83 1.89 0.83 1.89 1.38 1.83 1.38 1.83 0.32 1.89 0.32 1.89 0.77 1.95 0.77 ;
      POLYGON 1.685 1.38 1.625 1.38 1.625 0.585 1.12 0.585 1.12 1.165 1.24 1.165 1.24 1.38 0.905 1.38 0.905 1.165 1.06 1.165 1.06 0.585 0.725 0.585 0.725 0.595 0.695 0.595 0.695 1.035 0.725 1.035 0.725 1.095 0.605 1.095 0.605 1.035 0.635 1.035 0.635 0.595 0.605 0.595 0.605 0.535 0.635 0.535 0.635 0.525 1.185 0.525 1.185 0.32 1.245 0.32 1.245 0.525 1.625 0.525 1.625 0.32 1.685 0.32 ;
      POLYGON 1.335 0.705 1.305 0.705 1.305 1.035 1.335 1.035 1.335 1.095 1.215 1.095 1.215 1.035 1.245 1.035 1.245 0.705 1.215 0.705 1.215 0.645 1.335 0.645 ;
      POLYGON 1.32 3.115 1.26 3.115 1.26 2.6 0.98 2.6 0.98 2.54 1.26 2.54 1.26 2.185 1.32 2.185 ;
      POLYGON 0.93 1.095 0.81 1.095 0.81 1.035 0.84 1.035 0.84 0.72 0.9 0.72 0.9 1.035 0.93 1.035 ;
      POLYGON 0.91 3.115 0.85 3.115 0.85 2.625 0.79 2.625 0.79 2.505 0.85 2.505 0.85 2.185 0.91 2.185 ;
      POLYGON 0.64 2.1 0.57 2.1 0.57 3.115 0.51 3.115 0.51 2.015 0.61 2.015 0.61 2.04 0.64 2.04 ;
      POLYGON 0.45 1.52 0.29 1.52 0.29 1.46 0.39 1.46 0.39 0.32 0.45 0.32 ;
      RECT 0.1 0.135 0.16 1.2 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RDFFSQX1

MACRO RDFFSRQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RDFFSRQX1 0 0 ;
  SIZE 6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 1.77 5.73 1.77 5.73 2.46 5.67 2.46 5.67 1.77 1.56 1.77 1.56 2.385 1.5 2.385 1.5 1.77 1.115 1.77 1.115 2.4 1.055 2.4 1.055 1.77 0.26 1.77 0.26 2.4 0.2 2.4 0.2 1.77 -0.005 1.77 -0.005 1.65 0.89 1.65 0.89 1.27 0.95 1.27 0.95 1.65 1.68 1.65 1.68 1.27 1.74 1.27 1.74 1.65 5.23 1.65 5.23 1.13 5.29 1.13 5.29 1.65 5.745 1.65 5.745 1.13 5.805 1.13 5.805 1.65 6 1.65 ;
    END
  END VDD
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0516 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.5925925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 23.287037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.165 0.92 1.09 0.92 1.09 1.14 1.12 1.14 1.12 1.2 1 1.2 1 1.14 1.03 1.14 1.03 0.72 1.165 0.72 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.83333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.025 2.69 1.185 2.845 ;
    END
  END CK
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.695 2.61 3.215 2.61 3.215 2 3.345 2 3.345 1.89 3.595 1.89 3.595 2 3.695 2 ;
    END
  END ExtVDD
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.9074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.64 2.59 1.565 2.59 1.565 2.83 1.435 2.83 1.435 2.5 1.565 2.5 1.565 2.53 1.64 2.53 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.027225 LAYER Metal1 ;
    ANTENNADIFFAREA 3.6339 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.23985 LAYER Metal1 ;
      ANTENNAMAXAREACAR 20.95987075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 153.3208255 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.565 2.82 5.525 2.82 5.525 3.135 5.465 3.135 5.465 2.82 5.435 2.82 5.435 2.5 5.465 2.5 5.465 2.07 5.525 2.07 5.525 2.5 5.565 2.5 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.16 2.69 0.365 2.82 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 3.48 0 3.48 0 3.36 0.2 3.36 0.2 2.97 0.26 2.97 0.26 3.36 1.055 3.36 1.055 2.97 1.115 2.97 1.115 3.36 1.5 3.36 1.5 2.97 1.56 2.97 1.56 3.36 3.215 3.36 3.215 3.025 3.275 3.025 3.275 3.36 3.635 3.36 3.635 3.025 3.695 3.025 3.695 3.36 5.67 3.36 5.67 2.875 5.73 2.875 5.73 3.36 6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6 0.06 5.865 0.06 5.865 0.465 5.805 0.465 5.805 0.06 3.79 0.06 3.79 0.465 3.73 0.465 3.73 0.06 0.95 0.06 0.95 0.32 1.125 0.32 1.125 0.465 0.89 0.465 0.89 0.06 0 0.06 0 -0.06 6 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.10185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.41 1.525 4.255 1.525 4.255 1.37 4.11 1.37 4.11 0.41 4.17 0.41 4.17 1.31 4.41 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.66 0.465 5.6 0.465 5.6 0.26 5.25 0.26 5.25 0.465 5.19 0.465 5.19 0.2 5.66 0.2 ;
      POLYGON 5.6 1.345 5.54 1.345 5.54 1.015 5.05 1.015 5.05 1.345 4.99 1.345 4.99 0.955 5.6 0.955 ;
      POLYGON 5.455 0.67 4.99 0.67 4.99 0.32 5.05 0.32 5.05 0.61 5.395 0.61 5.395 0.32 5.455 0.32 ;
      RECT 4.785 0.32 4.845 1.345 ;
      RECT 4.095 2.385 4.54 2.445 ;
      POLYGON 4.535 1.13 4.265 1.13 4.265 0.25 4.255 0.25 4.255 0.23 4.24 0.23 4.24 0.17 4.255 0.17 4.255 0.13 4.315 0.13 4.315 0.17 4.325 0.17 4.325 1.07 4.535 1.07 ;
      RECT 4.445 0.135 4.505 0.995 ;
      POLYGON 4.195 1.51 3.935 1.51 3.935 0.83 3.4 0.83 3.4 0.245 3.46 0.245 3.46 0.77 3.935 0.77 3.935 0.32 3.995 0.32 3.995 1.45 4.195 1.45 ;
      POLYGON 4.005 3.17 3.945 3.17 3.945 2.78 3.145 2.78 3.145 2.72 3.945 2.72 3.945 2 4.005 2 ;
      POLYGON 3.8 2.93 3.07 2.93 3.07 3.17 3.01 3.17 3.01 2 3.07 2 3.07 2.87 3.8 2.87 ;
      RECT 3.51 1.24 3.79 1.525 ;
      RECT 3.215 0.32 3.275 1.455 ;
      POLYGON 3.07 1.52 2.78 1.52 2.78 1.46 3.01 1.46 3.01 0.32 3.07 0.32 ;
      RECT 2.475 0.6 2.535 1.285 ;
      POLYGON 2.245 0.83 2.185 0.83 2.185 1.485 2.125 1.485 2.125 0.32 2.185 0.32 2.185 0.77 2.245 0.77 ;
      POLYGON 2.065 1.19 1.98 1.19 1.98 1.485 1.92 1.485 1.92 1.13 2.005 1.13 2.005 0.585 1.31 0.585 1.31 1.27 1.43 1.27 1.43 1.485 1.095 1.485 1.095 1.27 1.25 1.27 1.25 0.585 0.915 0.585 0.915 0.595 0.885 0.595 0.885 1.14 0.915 1.14 0.915 1.2 0.795 1.2 0.795 1.14 0.825 1.14 0.825 0.595 0.795 0.595 0.795 0.535 0.825 0.535 0.825 0.525 1.475 0.525 1.475 0.32 1.535 0.32 1.535 0.525 1.92 0.525 1.92 0.32 1.98 0.32 1.98 0.525 2.065 0.525 ;
      POLYGON 1.915 0.705 1.875 0.705 1.875 0.75 1.86 0.75 1.86 1.18 1.8 1.18 1.8 0.705 1.795 0.705 1.795 0.645 1.915 0.645 ;
      POLYGON 1.805 2.57 1.765 2.57 1.765 3.115 1.705 3.115 1.705 2.17 1.765 2.17 1.765 2.45 1.805 2.45 ;
      POLYGON 1.775 0.465 1.715 0.465 1.715 0.255 1.33 0.255 1.33 0.465 1.27 0.465 1.27 0.195 1.775 0.195 ;
      POLYGON 1.715 0.705 1.685 0.705 1.685 1.185 1.525 1.185 1.525 1.2 1.405 1.2 1.405 1.14 1.435 1.14 1.435 1.125 1.625 1.125 1.625 0.705 1.595 0.705 1.595 0.645 1.715 0.645 ;
      POLYGON 1.32 3.115 1.26 3.115 1.26 2.6 0.98 2.6 0.98 2.54 1.26 2.54 1.26 2.185 1.32 2.185 ;
      POLYGON 0.91 3.115 0.85 3.115 0.85 2.625 0.79 2.625 0.79 2.505 0.85 2.505 0.85 2.185 0.91 2.185 ;
      POLYGON 0.64 1.525 0.37 1.525 0.37 1.465 0.58 1.465 0.58 0.32 0.64 0.32 ;
      POLYGON 0.64 2.075 0.57 2.075 0.57 3.115 0.51 3.115 0.51 2.015 0.64 2.015 ;
      RECT 0.28 0.135 0.34 1.305 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RDFFSRQX1

MACRO RDFFSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RDFFSRX1 0 0 ;
  SIZE 6.2 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 5.935 1.77 5.935 2.46 5.875 2.46 5.875 1.77 5.255 1.77 5.255 2.46 5.195 2.46 5.195 1.77 1.465 1.77 1.465 2.28 1.405 2.28 1.405 1.77 0.62 1.77 0.62 2.28 0.56 2.28 0.56 1.77 0 1.77 0 1.65 0.25 1.65 0.25 1.05 0.31 1.05 0.31 1.65 1.095 1.65 1.095 1.27 1.155 1.27 1.155 1.65 1.25 1.65 1.25 1.27 1.31 1.27 1.31 1.65 1.885 1.65 1.885 1.27 1.945 1.27 1.945 1.65 5.435 1.65 5.435 1.13 5.495 1.13 5.495 1.65 5.95 1.65 5.95 1.13 6.01 1.13 6.01 1.65 6.2 1.65 ;
    END
  END VDD
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.116 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 3.580247 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 36.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 0.92 1.31 0.92 1.31 1.14 1.34 1.14 1.34 1.2 1.22 1.2 1.22 1.14 1.25 1.14 1.25 0.92 1.235 0.92 1.235 0.72 1.365 0.72 ;
    END
  END SN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 3.42 2 3.9 2.61 ;
    END
  END ExtVDD
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.85185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.39 0.905 0.38 0.905 0.38 0.98 0.26 0.98 0.26 0.74 0.38 0.74 0.38 0.845 0.39 0.845 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6253 LAYER Metal1 ;
    ANTENNADIFFAREA 3.76965 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2853 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.71713975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 151.77707675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.765 2.82 5.73 2.82 5.73 3.135 5.67 3.135 5.67 2.82 5.635 2.82 5.635 2.69 5.67 2.69 5.67 2.07 5.73 2.07 5.73 2.69 5.765 2.69 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6253 LAYER Metal1 ;
    ANTENNADIFFAREA 3.76965 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2853 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.71713975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 151.77707675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.05 3.135 4.99 3.135 4.99 2.63 4.835 2.63 4.835 2.5 4.99 2.5 4.99 2.07 5.05 2.07 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.31481475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 2.66 0.67 2.82 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 3.48 0 3.48 0 3.36 0.56 3.36 0.56 2.97 0.62 2.97 0.62 3.36 1.405 3.36 1.405 2.97 1.465 2.97 1.465 3.36 3.42 3.36 3.42 3.025 3.48 3.025 3.48 3.36 3.84 3.36 3.84 3.025 3.9 3.025 3.9 3.36 5.195 3.36 5.195 2.875 5.255 2.875 5.255 3.36 5.875 3.36 5.875 2.875 5.935 2.875 5.935 3.36 6.2 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 6.07 0.06 6.07 0.465 6.01 0.465 6.01 0.06 3.955 0.06 3.955 0.34 3.895 0.34 3.895 0.06 1.155 0.06 1.155 0.32 1.33 0.32 1.33 0.465 1.095 0.465 1.095 0.06 0.31 0.06 0.31 0.465 0.25 0.465 0.25 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.29629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.405 2.69 1.565 2.87 ;
    END
  END CK
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.62962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.46 1.095 4.755 1.3 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.865 0.465 5.805 0.465 5.805 0.26 5.455 0.26 5.455 0.465 5.395 0.465 5.395 0.2 5.865 0.2 ;
      POLYGON 5.805 1.345 5.745 1.345 5.745 1.015 5.255 1.015 5.255 1.345 5.195 1.345 5.195 0.955 5.805 0.955 ;
      POLYGON 5.66 0.67 5.195 0.67 5.195 0.32 5.255 0.32 5.255 0.61 5.6 0.61 5.6 0.32 5.66 0.32 ;
      POLYGON 5.49 3.075 5.43 3.075 5.43 2.685 5.135 2.685 5.135 2.625 5.43 2.625 5.43 2.155 5.49 2.155 ;
      POLYGON 5.05 1.345 4.99 1.345 4.99 0.425 4.775 0.425 4.775 0.365 4.99 0.365 4.99 0.32 5.05 0.32 ;
      POLYGON 5.025 1.55 2.61 1.55 2.61 1.025 2.67 1.025 2.67 1.49 5.025 1.49 ;
      POLYGON 4.905 0.665 4.875 0.665 4.875 1.425 2.78 1.425 2.78 1.365 4.815 1.365 4.815 0.665 4.785 0.665 4.785 0.605 4.815 0.605 4.815 0.51 4.875 0.51 4.875 0.605 4.905 0.605 ;
      RECT 4.3 2.385 4.745 2.445 ;
      POLYGON 4.715 1 4.47 1 4.47 0.25 4.46 0.25 4.46 0.23 4.445 0.23 4.445 0.17 4.46 0.17 4.46 0.13 4.52 0.13 4.52 0.17 4.53 0.17 4.53 0.94 4.715 0.94 ;
      RECT 4.65 0.135 4.71 0.84 ;
      POLYGON 4.37 1.235 4.31 1.235 4.31 1.22 4.2 1.22 4.2 1.255 4.14 1.255 4.14 1.13 4.2 1.13 4.2 1.16 4.31 1.16 4.31 0.415 4.2 0.415 4.2 0.47 3.715 0.47 3.715 0.3 3.6 0.3 3.6 0.24 3.775 0.24 3.775 0.41 4.14 0.41 4.14 0.32 4.2 0.32 4.2 0.355 4.37 0.355 ;
      POLYGON 4.245 0.68 4.185 0.68 4.185 0.65 3.615 0.65 3.615 0.59 4.185 0.59 4.185 0.56 4.245 0.56 ;
      POLYGON 4.245 0.89 4.185 0.89 4.185 0.86 3.85 0.86 3.85 0.8 4.185 0.8 4.185 0.77 4.245 0.77 ;
      POLYGON 4.21 3.17 4.15 3.17 4.15 2.78 3.35 2.78 3.35 2.72 4.15 2.72 4.15 2 4.21 2 ;
      POLYGON 4.005 2.93 3.275 2.93 3.275 3.17 3.215 3.17 3.215 2 3.275 2 3.275 2.87 4.005 2.87 ;
      RECT 3.74 1.13 3.995 1.25 ;
      POLYGON 3.655 1.25 3.42 1.25 3.42 0.32 3.48 0.32 3.48 1.19 3.595 1.19 3.595 1.13 3.655 1.13 ;
      POLYGON 3.275 1.255 3.215 1.255 3.215 0.65 2.39 0.65 2.39 1.485 2.33 1.485 2.33 0.32 2.39 0.32 2.39 0.59 3.155 0.59 3.155 0.58 3.215 0.58 3.215 0.32 3.275 0.32 ;
      POLYGON 2.27 1.19 2.185 1.19 2.185 1.485 2.125 1.485 2.125 1.13 2.21 1.13 2.21 0.585 1.515 0.585 1.515 1.27 1.635 1.27 1.635 1.485 1.455 1.485 1.455 0.585 1.12 0.585 1.12 0.595 1.09 0.595 1.09 1.14 1.12 1.14 1.12 1.2 1 1.2 1 1.14 1.03 1.14 1.03 0.595 1 0.595 1 0.535 1.03 0.535 1.03 0.525 1.68 0.525 1.68 0.32 1.74 0.32 1.74 0.525 2.125 0.525 2.125 0.32 2.185 0.32 2.185 0.525 2.27 0.525 ;
      POLYGON 2.12 0.705 2.08 0.705 2.08 0.75 2.065 0.75 2.065 1.18 2.005 1.18 2.005 0.705 2 0.705 2 0.645 2.12 0.645 ;
      POLYGON 1.98 0.465 1.92 0.465 1.92 0.255 1.535 0.255 1.535 0.465 1.475 0.465 1.475 0.195 1.98 0.195 ;
      POLYGON 1.92 0.705 1.89 0.705 1.89 1.185 1.61 1.185 1.61 1.125 1.83 1.125 1.83 0.705 1.8 0.705 1.8 0.645 1.92 0.645 ;
      POLYGON 1.73 3.03 1.67 3.03 1.67 3.115 1.61 3.115 1.61 2.97 1.67 2.97 1.67 2.565 1.33 2.565 1.33 2.505 1.67 2.505 1.67 2.28 1.61 2.28 1.61 2.065 1.67 2.065 1.67 2.13 1.73 2.13 ;
      POLYGON 1.26 3.115 1.2 3.115 1.2 2.66 1.14 2.66 1.14 2.54 1.2 2.54 1.2 2.065 1.26 2.065 ;
      POLYGON 0.93 3.115 0.87 3.115 0.87 2.435 0.345 2.435 0.345 2.375 0.87 2.375 0.87 2.065 0.93 2.065 ;
      POLYGON 0.845 1.485 0.435 1.485 0.435 1.56 0.375 1.56 0.375 1.425 0.785 1.425 0.785 0.32 0.845 0.32 ;
      RECT 0.615 0.135 0.675 1.305 ;
      POLYGON 0.555 0.985 0.515 0.985 0.515 1.265 0.455 1.265 0.455 0.32 0.515 0.32 0.515 0.865 0.555 0.865 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RDFFSRX1

MACRO RDFFSX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RDFFSX1 0 0 ;
  SIZE 5.8 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 1.77 5.53 1.77 5.53 2.46 5.47 2.46 5.47 1.77 4.85 1.77 4.85 2.46 4.79 2.46 4.79 1.77 1.115 1.77 1.115 2.4 1.055 2.4 1.055 1.77 0.26 1.77 0.26 2.4 0.2 2.4 0.2 1.77 -0.005 1.77 -0.005 1.65 0.7 1.65 0.7 1.165 0.76 1.165 0.76 1.65 1.38 1.65 1.38 1.25 1.385 1.25 1.385 1.165 1.445 1.165 1.445 1.38 1.44 1.38 1.44 1.65 5.03 1.65 5.03 1.13 5.09 1.13 5.09 1.65 5.44 1.65 5.44 1.13 5.5 1.13 5.5 1.65 5.8 1.65 ;
    END
  END VDD
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0516 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.5925925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 21.9444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.965 1.095 0.81 1.095 0.81 1.035 0.82 1.035 0.82 0.79 0.84 0.79 0.84 0.72 0.9 0.72 0.9 0.79 0.965 0.79 ;
    END
  END SN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.495 2.61 3.015 2.61 3.015 2 3.145 2 3.145 1.89 3.395 1.89 3.395 2 3.495 2 ;
    END
  END ExtVDD
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.64814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.035 2.69 1.185 2.845 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.80595 LAYER Metal1 ;
    ANTENNADIFFAREA 3.6343 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2529 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.003361 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 137.995255 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.365 2.82 5.325 2.82 5.325 3.135 5.265 3.135 5.265 2.82 5.235 2.82 5.235 2.69 5.265 2.69 5.265 2.07 5.325 2.07 5.325 2.69 5.365 2.69 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.80595 LAYER Metal1 ;
    ANTENNADIFFAREA 3.6343 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2529 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.003361 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 137.995255 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.645 3.135 4.585 3.135 4.585 2.63 4.435 2.63 4.435 2.5 4.585 2.5 4.585 2.07 4.645 2.07 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.462963 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.2 2.69 0.365 2.82 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 3.48 0 3.48 0 3.36 0.2 3.36 0.2 2.97 0.26 2.97 0.26 3.36 1.055 3.36 1.055 2.97 1.115 2.97 1.115 3.36 3.015 3.36 3.015 3.025 3.075 3.025 3.075 3.36 3.435 3.36 3.435 3.025 3.495 3.025 3.495 3.36 4.79 3.36 4.79 2.875 4.85 2.875 4.85 3.36 5.47 3.36 5.47 2.875 5.53 2.875 5.53 3.36 5.8 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 0.06 5.5 0.06 5.5 0.465 5.44 0.465 5.44 0.06 3.59 0.06 3.59 0.465 3.53 0.465 3.53 0.06 0.76 0.06 0.76 0.32 0.935 0.32 0.935 0.465 0.7 0.465 0.7 0.06 0 0.06 0 -0.06 5.8 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.7685185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.39 1.525 4.055 1.525 4.055 1.37 3.91 1.37 3.91 0.41 3.97 0.41 3.97 1.31 4.39 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.295 1.345 5.235 1.345 5.235 1.015 4.85 1.015 4.85 1.345 4.79 1.345 4.79 0.955 5.295 0.955 ;
      POLYGON 5.19 0.465 5.13 0.465 5.13 0.42 4.85 0.42 4.85 0.495 4.79 0.495 4.79 0.32 4.85 0.32 4.85 0.36 5.13 0.36 5.13 0.32 5.19 0.32 ;
      POLYGON 5.085 3.08 5.025 3.08 5.025 2.655 4.73 2.655 4.73 2.595 5.025 2.595 5.025 2.16 5.085 2.16 ;
      RECT 4.585 0.32 4.645 1.345 ;
      RECT 3.895 2.385 4.34 2.445 ;
      POLYGON 4.335 1.13 4.065 1.13 4.065 0.25 4.055 0.25 4.055 0.23 4.04 0.23 4.04 0.17 4.055 0.17 4.055 0.13 4.115 0.13 4.115 0.17 4.125 0.17 4.125 1.07 4.335 1.07 ;
      RECT 4.245 0.135 4.305 0.995 ;
      POLYGON 3.995 1.51 3.735 1.51 3.735 0.83 3.2 0.83 3.2 0.245 3.26 0.245 3.26 0.77 3.735 0.77 3.735 0.32 3.795 0.32 3.795 1.45 3.995 1.45 ;
      POLYGON 3.805 3.17 3.745 3.17 3.745 2.78 2.945 2.78 2.945 2.72 3.745 2.72 3.745 2 3.805 2 ;
      POLYGON 3.6 2.93 2.87 2.93 2.87 3.17 2.81 3.17 2.81 2 2.87 2 2.87 2.87 3.6 2.87 ;
      RECT 3.31 1.24 3.59 1.525 ;
      RECT 3.015 0.32 3.075 1.455 ;
      POLYGON 2.87 1.52 2.58 1.52 2.58 1.46 2.81 1.46 2.81 0.32 2.87 0.32 ;
      RECT 2.275 0.6 2.335 1.18 ;
      POLYGON 1.95 0.83 1.89 0.83 1.89 1.38 1.83 1.38 1.83 0.32 1.89 0.32 1.89 0.77 1.95 0.77 ;
      POLYGON 1.685 1.38 1.625 1.38 1.625 0.585 1.12 0.585 1.12 1.165 1.24 1.165 1.24 1.38 0.905 1.38 0.905 1.165 1.06 1.165 1.06 0.585 0.725 0.585 0.725 0.595 0.695 0.595 0.695 1.035 0.725 1.035 0.725 1.095 0.605 1.095 0.605 1.035 0.635 1.035 0.635 0.595 0.605 0.595 0.605 0.535 0.635 0.535 0.635 0.525 1.185 0.525 1.185 0.32 1.245 0.32 1.245 0.525 1.625 0.525 1.625 0.32 1.685 0.32 ;
      POLYGON 1.335 0.705 1.305 0.705 1.305 1.035 1.335 1.035 1.335 1.095 1.215 1.095 1.215 1.035 1.245 1.035 1.245 0.705 1.215 0.705 1.215 0.645 1.335 0.645 ;
      POLYGON 1.32 3.115 1.26 3.115 1.26 2.6 0.98 2.6 0.98 2.54 1.26 2.54 1.26 2.185 1.32 2.185 ;
      POLYGON 0.91 3.115 0.85 3.115 0.85 2.63 0.79 2.63 0.79 2.51 0.85 2.51 0.85 2.185 0.91 2.185 ;
      POLYGON 0.64 2.1 0.57 2.1 0.57 3.115 0.51 3.115 0.51 2.015 0.61 2.015 0.61 2.04 0.64 2.04 ;
      POLYGON 0.45 1.52 0.29 1.52 0.29 1.46 0.39 1.46 0.39 0.32 0.45 0.32 ;
      RECT 0.1 0.135 0.16 1.2 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RDFFSX1

MACRO RDFFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RDFFX1 0 0 ;
  SIZE 5.2 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.2 1.77 4.93 1.77 4.93 2.46 4.87 2.46 4.87 1.77 4.255 1.77 4.255 2.465 4.195 2.465 4.195 1.77 1.035 1.77 1.035 2.4 0.975 2.4 0.975 1.77 0.255 1.77 0.255 2.4 0.195 2.4 0.195 1.77 0 1.77 0 1.65 0.895 1.65 0.895 1.11 0.955 1.11 0.955 1.65 4.3 1.65 4.3 1.13 4.36 1.13 4.36 1.65 5.2 1.65 ;
    END
  END VDD
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2354 LAYER Metal1 ;
    ANTENNADIFFAREA 3.206275 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2529 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.747331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 121.376038 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.05 3.13 3.99 3.13 3.99 2.63 3.835 2.63 3.835 2.5 3.99 2.5 3.99 2.075 4.05 2.075 ;
    END
  END QN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.9 2.61 2.42 2.61 2.42 2 2.57 2 2.57 1.89 2.82 1.89 2.82 2 2.9 2 ;
    END
  END ExtVDD
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2354 LAYER Metal1 ;
    ANTENNADIFFAREA 3.206275 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2529 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.747331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 121.376038 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.765 2.82 4.725 2.82 4.725 3.135 4.665 3.135 4.665 2.82 4.635 2.82 4.635 2.69 4.665 2.69 4.665 2.07 4.725 2.07 4.725 2.69 4.765 2.69 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.4814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.185 2.65 0.365 2.82 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.2 3.48 0 3.48 0 3.36 0.195 3.36 0.195 2.97 0.255 2.97 0.255 3.36 0.975 3.36 0.975 2.97 1.035 2.97 1.035 3.36 2.42 3.36 2.42 3.025 2.48 3.025 2.48 3.36 2.84 3.36 2.84 3.025 2.9 3.025 2.9 3.36 4.195 3.36 4.195 2.87 4.255 2.87 4.255 3.36 4.87 3.36 4.87 2.875 4.93 2.875 4.93 3.36 5.2 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.2 0.06 4.36 0.06 4.36 0.465 4.3 0.465 4.3 0.06 2.995 0.06 2.995 0.625 2.935 0.625 2.935 0.06 0.955 0.06 0.955 0.54 0.895 0.54 0.895 0.06 0 0.06 0 -0.06 5.2 -0.06 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.985 2.5 1.165 2.645 ;
    END
  END CK
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0933 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.87962975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 22.962963 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.46 1.155 3.7 1.36 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 4.49 3.075 4.43 3.075 4.43 2.685 4.135 2.685 4.135 2.625 4.43 2.625 4.43 2.165 4.49 2.165 ;
      POLYGON 4.05 1.345 3.99 1.345 3.99 1.05 3.96 1.05 3.96 0.93 3.99 0.93 3.99 0.32 4.05 0.32 ;
      RECT 3.775 0.14 3.835 1.45 ;
      RECT 3.3 2.615 3.745 2.675 ;
      POLYGON 3.42 1.525 3.14 1.525 3.14 1.025 2.66 1.025 2.66 0.38 2.72 0.38 2.72 0.965 3.14 0.965 3.14 0.48 3.2 0.48 3.2 1.465 3.42 1.465 ;
      RECT 3.31 0.48 3.37 1.215 ;
      POLYGON 3.21 3.17 3.15 3.17 3.15 2.78 2.35 2.78 2.35 2.72 3.15 2.72 3.15 2 3.21 2 ;
      POLYGON 3.005 2.93 2.275 2.93 2.275 3.17 2.215 3.17 2.215 2 2.275 2 2.275 2.87 3.005 2.87 ;
      POLYGON 2.995 1.555 2.735 1.555 2.735 1.26 2.935 1.26 2.935 1.255 2.995 1.255 ;
      RECT 2.42 0.48 2.48 1.47 ;
      POLYGON 2.275 1.54 2.005 1.54 2.005 1.48 2.215 1.48 2.215 0.48 2.275 0.48 ;
      POLYGON 2.125 1.02 2.005 1.02 2.005 0.96 2.035 0.96 2.035 0.86 1.365 0.86 1.365 1.325 1.305 1.325 1.305 0.38 1.365 0.38 1.365 0.8 2.095 0.8 2.095 0.96 2.125 0.96 ;
      POLYGON 1.3 3.03 1.24 3.03 1.24 3.115 1.18 3.115 1.18 2.97 1.24 2.97 1.24 2.795 0.895 2.795 0.895 2.735 1.24 2.735 1.24 2.4 1.18 2.4 1.18 2.185 1.24 2.185 1.24 2.25 1.3 2.25 ;
      POLYGON 1.16 1.325 1.1 1.325 1.1 0.85 0.89 0.85 0.89 0.98 0.92 0.98 0.92 1.04 0.8 1.04 0.8 0.98 0.83 0.98 0.83 0.67 0.8 0.67 0.8 0.61 0.92 0.61 0.92 0.67 0.89 0.67 0.89 0.79 1.1 0.79 1.1 0.395 1.16 0.395 ;
      POLYGON 0.83 3.115 0.77 3.115 0.77 2.62 0.68 2.62 0.68 2.56 0.77 2.56 0.77 2.185 0.83 2.185 ;
      POLYGON 0.645 1.325 0.635 1.325 0.635 1.525 0.475 1.525 0.475 1.465 0.575 1.465 0.575 1.11 0.585 1.11 0.585 0.395 0.645 0.395 ;
      POLYGON 0.61 2.155 0.565 2.155 0.565 3.115 0.505 3.115 0.505 2.095 0.55 2.095 0.55 1.84 0.61 1.84 ;
      RECT 0.305 0.145 0.365 1.545 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RDFFX1

MACRO RTLATRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RTLATRX1 0 0 ;
  SIZE 5 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.755 2.61 2.56 2.61 2.56 2.635 2.43 2.635 2.43 2.61 2.225 2.61 2.225 1.92 2.38 1.92 2.38 1.98 2.285 1.98 2.285 2.31 2.695 2.31 2.695 2.125 2.755 2.125 ;
    END
  END ExtVDD
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 1.77 4.665 1.77 4.665 2.46 4.605 2.46 4.605 1.77 4.2 1.77 4.2 2.46 4.14 2.46 4.14 1.77 0.43 1.77 0.43 2.27 0.37 2.27 0.37 1.77 0 1.77 0 1.65 0.425 1.65 0.425 1.17 0.485 1.17 0.485 1.65 4.405 1.65 4.405 1.15 4.465 1.15 4.465 1.65 4.815 1.65 4.815 1.15 4.875 1.15 4.875 1.65 5 1.65 ;
    END
  END VDD
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.7314815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.22 0.595 0.38 0.73 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.91875 LAYER Metal1 ;
    ANTENNADIFFAREA 2.8113 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20115 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.48173 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 147.56152125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.93 2.885 4.87 2.885 4.87 3.155 4.81 3.155 4.81 2.825 4.87 2.825 4.87 2.65 4.81 2.65 4.81 2.07 4.87 2.07 4.87 2.59 4.93 2.59 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.91875 LAYER Metal1 ;
    ANTENNADIFFAREA 2.791 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20115 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.48173 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 147.56152125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.995 3.155 3.935 3.155 3.935 3.01 3.835 3.01 3.835 2.69 3.935 2.69 3.935 2.07 3.995 2.07 ;
    END
  END QN
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.462963 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.79 0.58 0.94 ;
    END
  END G
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.42 2.495 0.575 2.63 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 3.48 0 3.48 0 3.36 0.37 3.36 0.37 2.975 0.43 2.975 0.43 3.36 1.92 3.36 1.92 2.95 1.98 2.95 1.98 3.36 2.895 3.36 2.895 2.89 2.955 2.89 2.955 3.36 4.14 3.36 4.14 2.895 4.2 2.895 4.2 3.36 4.605 3.36 4.605 2.895 4.665 2.895 4.665 3.36 5 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5 0.06 4.875 0.06 4.875 0.545 4.815 0.545 4.815 0.06 2.54 0.06 2.54 0.49 2.48 0.49 2.48 0.06 0.28 0.06 0.28 0.495 0.22 0.495 0.22 0.06 0 0.06 0 -0.06 5 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0942 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.9074075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 33.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 0.97 1.655 1.11 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 4.67 1.365 4.61 1.365 4.61 1.055 4.21 1.055 4.21 1.365 4.15 1.365 4.15 0.995 4.67 0.995 ;
      POLYGON 4.565 0.64 4.245 0.64 4.245 0.4 4.305 0.4 4.305 0.58 4.505 0.58 4.505 0.4 4.565 0.4 ;
      POLYGON 4.495 2.755 4.405 2.755 4.405 3.155 4.345 3.155 4.345 2.07 4.405 2.07 4.405 2.695 4.495 2.695 ;
      POLYGON 4.1 0.905 4.005 0.905 4.005 1.365 3.945 1.365 3.945 0.905 2.37 0.905 2.37 0.845 4.04 0.845 4.04 0.4 4.1 0.4 ;
      RECT 1.445 1.485 3.71 1.545 ;
      RECT 2.155 0.7 3.31 0.76 ;
      POLYGON 3.215 2.87 3.155 2.87 3.155 1.96 2.555 1.96 2.555 1.9 3.215 1.9 ;
      POLYGON 3.065 2.82 2.645 2.82 2.645 3.035 2.585 3.035 2.585 2.875 2.37 2.875 2.37 2.815 2.585 2.815 2.585 2.76 3.005 2.76 3.005 2.125 3.065 2.125 ;
      POLYGON 2.995 0.61 2.25 0.61 2.25 0.49 2.31 0.49 2.31 0.55 2.685 0.55 2.685 0.345 2.745 0.345 2.745 0.55 2.995 0.55 ;
      POLYGON 2.995 1.23 2.745 1.23 2.745 1.305 2.685 1.305 2.685 1.09 2.745 1.09 2.745 1.17 2.995 1.17 ;
      POLYGON 2.54 1.395 2.375 1.395 2.375 1.42 2.315 1.42 2.315 1.3 2.375 1.3 2.375 1.335 2.48 1.335 2.48 1.09 2.54 1.09 ;
      POLYGON 2.29 1.2 2.08 1.2 2.08 1.305 2.02 1.305 2.02 0.355 2.08 0.355 2.08 1.14 2.29 1.14 ;
      POLYGON 2.265 2.73 2.185 2.73 2.185 3.095 2.125 3.095 2.125 2.73 2.02 2.73 2.02 2.125 2.08 2.125 2.08 2.67 2.265 2.67 ;
      POLYGON 1.875 1.335 1.05 1.335 1.05 1.275 1.815 1.275 1.815 0.355 1.875 0.355 ;
      POLYGON 1.17 2.385 0.84 2.385 0.84 3.035 0.74 3.035 0.74 3.12 0.68 3.12 0.68 2.975 0.78 2.975 0.78 2.385 0.68 2.385 0.68 2.055 0.74 2.055 0.74 2.325 1.17 2.325 ;
      POLYGON 0.87 0.76 0.75 0.76 0.75 1.23 0.69 1.23 0.69 1.385 0.63 1.385 0.63 1.17 0.69 1.17 0.69 1.1 0.28 1.1 0.28 1.545 0.09 1.545 0.09 1.485 0.22 1.485 0.22 1.04 0.69 1.04 0.69 0.58 0.53 0.58 0.53 0.35 0.59 0.35 0.59 0.52 0.75 0.52 0.75 0.7 0.87 0.7 ;
      POLYGON 0.695 2.845 0.225 2.845 0.225 3.12 0.165 3.12 0.165 2.055 0.225 2.055 0.225 2.785 0.695 2.785 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RTLATRX1

MACRO RTLATSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RTLATSRX1 0 0 ;
  SIZE 5 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.765 2.63 2.435 2.63 2.435 2.61 2.225 2.61 2.225 1.98 1.875 1.98 1.875 2.34 1.815 2.34 1.815 1.92 2.38 1.92 2.38 1.98 2.285 1.98 2.285 2.31 2.695 2.31 2.695 2.125 2.755 2.125 2.755 2.31 2.765 2.31 ;
    END
  END ExtVDD
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 1.77 4.665 1.77 4.665 2.46 4.605 2.46 4.605 1.77 4.2 1.77 4.2 2.46 4.14 2.46 4.14 1.77 0.43 1.77 0.43 2.27 0.37 2.27 0.37 1.77 0 1.77 0 1.65 0.425 1.65 0.425 1.17 0.485 1.17 0.485 1.65 4.405 1.65 4.405 1.15 4.465 1.15 4.465 1.65 4.815 1.65 4.815 1.15 4.875 1.15 4.875 1.65 5 1.65 ;
    END
  END VDD
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.824074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.22 0.58 0.375 0.73 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.976775 LAYER Metal1 ;
    ANTENNADIFFAREA 2.8544 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20115 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.77019625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 149.9627145 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.93 2.87 4.87 2.87 4.87 3.155 4.81 3.155 4.81 2.81 4.87 2.81 4.87 2.65 4.81 2.65 4.81 2.07 4.87 2.07 4.87 2.59 4.93 2.59 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.976775 LAYER Metal1 ;
    ANTENNADIFFAREA 2.8341 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20115 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.77019625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 149.9627145 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.995 3.155 3.935 3.155 3.935 3.01 3.835 3.01 3.835 2.69 3.935 2.69 3.935 2.07 3.995 2.07 ;
    END
  END QN
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.64814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.42 0.79 0.575 0.94 ;
    END
  END G
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.70370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.635 2.69 1.965 2.83 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.29629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.41 2.495 0.605 2.64 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 3.48 0 3.48 0 3.36 0.37 3.36 0.37 2.975 0.43 2.975 0.43 3.36 1.815 3.36 1.815 2.95 1.875 2.95 1.875 3.36 2.895 3.36 2.895 2.89 2.955 2.89 2.955 3.36 4.14 3.36 4.14 2.895 4.2 2.895 4.2 3.36 4.605 3.36 4.605 2.895 4.665 2.895 4.665 3.36 5 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5 0.06 4.875 0.06 4.875 0.545 4.815 0.545 4.815 0.06 2.54 0.06 2.54 0.49 2.48 0.49 2.48 0.06 0.28 0.06 0.28 0.495 0.22 0.495 0.22 0.06 0 0.06 0 -0.06 5 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0942 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.9074075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 33.70370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.415 0.97 1.655 1.11 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 4.67 1.365 4.61 1.365 4.61 1.055 4.21 1.055 4.21 1.365 4.15 1.365 4.15 0.995 4.67 0.995 ;
      POLYGON 4.565 0.64 4.245 0.64 4.245 0.4 4.305 0.4 4.305 0.58 4.505 0.58 4.505 0.4 4.565 0.4 ;
      POLYGON 4.495 2.755 4.405 2.755 4.405 3.155 4.345 3.155 4.345 2.07 4.405 2.07 4.405 2.695 4.495 2.695 ;
      POLYGON 4.1 0.905 4.005 0.905 4.005 1.365 3.945 1.365 3.945 0.905 2.37 0.905 2.37 0.845 4.04 0.845 4.04 0.4 4.1 0.4 ;
      RECT 1.445 1.485 3.71 1.545 ;
      RECT 2.155 0.7 3.31 0.76 ;
      POLYGON 3.215 2.87 3.155 2.87 3.155 1.96 2.555 1.96 2.555 1.9 3.215 1.9 ;
      POLYGON 3.065 2.82 2.645 2.82 2.645 3.035 2.585 3.035 2.585 2.875 2.37 2.875 2.37 2.815 2.585 2.815 2.585 2.76 3.005 2.76 3.005 2.125 3.065 2.125 ;
      POLYGON 2.995 0.61 2.25 0.61 2.25 0.49 2.31 0.49 2.31 0.55 2.685 0.55 2.685 0.345 2.745 0.345 2.745 0.55 2.995 0.55 ;
      POLYGON 2.995 1.23 2.745 1.23 2.745 1.305 2.685 1.305 2.685 1.09 2.745 1.09 2.745 1.17 2.995 1.17 ;
      POLYGON 2.54 1.395 2.375 1.395 2.375 1.42 2.315 1.42 2.315 1.3 2.375 1.3 2.375 1.335 2.48 1.335 2.48 1.09 2.54 1.09 ;
      POLYGON 2.29 1.2 2.08 1.2 2.08 1.305 2.02 1.305 2.02 0.355 2.08 0.355 2.08 1.14 2.29 1.14 ;
      POLYGON 2.28 2.73 2.14 2.73 2.14 2.95 2.185 2.95 2.185 3.095 2.125 3.095 2.125 3.04 2.08 3.04 2.08 2.495 2.02 2.495 2.02 2.125 2.08 2.125 2.08 2.435 2.15 2.435 2.15 2.495 2.14 2.495 2.14 2.67 2.28 2.67 ;
      POLYGON 1.875 1.335 1.05 1.335 1.05 1.275 1.815 1.275 1.815 0.355 1.875 0.355 ;
      POLYGON 1.17 2.385 0.84 2.385 0.84 3.035 0.74 3.035 0.74 3.12 0.68 3.12 0.68 2.975 0.78 2.975 0.78 2.385 0.68 2.385 0.68 2.055 0.74 2.055 0.74 2.325 1.17 2.325 ;
      POLYGON 0.92 0.76 0.705 0.76 0.705 1.385 0.63 1.385 0.63 1.17 0.645 1.17 0.645 1.1 0.28 1.1 0.28 1.545 0.09 1.545 0.09 1.485 0.22 1.485 0.22 1.04 0.645 1.04 0.645 0.495 0.53 0.495 0.53 0.35 0.59 0.35 0.59 0.435 0.705 0.435 0.705 0.7 0.92 0.7 ;
      POLYGON 0.695 2.845 0.225 2.845 0.225 3.12 0.165 3.12 0.165 2.055 0.225 2.055 0.225 2.785 0.695 2.785 ;
  END
  PROPERTY oaTaper "__DerivedDefaultTaperCG" ;
END RTLATSRX1

MACRO RTLATX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN RTLATX1 0 0 ;
  SIZE 5 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.765 2.63 2.415 2.63 2.415 2.61 2.225 2.61 2.225 1.92 2.38 1.92 2.38 1.98 2.285 1.98 2.285 2.31 2.695 2.31 2.695 2.125 2.755 2.125 2.755 2.31 2.765 2.31 ;
    END
  END ExtVDD
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 1.77 4.665 1.77 4.665 2.46 4.605 2.46 4.605 1.77 4.2 1.77 4.2 2.46 4.14 2.46 4.14 1.77 0.43 1.77 0.43 2.27 0.37 2.27 0.37 1.77 0 1.77 0 1.65 0.425 1.65 0.425 1.17 0.485 1.17 0.485 1.65 4.61 1.65 4.61 1.15 4.67 1.15 4.67 1.65 5 1.65 ;
    END
  END VDD
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6405 LAYER Metal1 ;
    ANTENNADIFFAREA 2.6459 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20115 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.098434 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 133.04996275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.93 2.88 4.87 2.88 4.87 3.155 4.81 3.155 4.81 2.82 4.87 2.82 4.87 2.69 4.81 2.69 4.81 2.07 4.87 2.07 4.87 2.63 4.93 2.63 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6405 LAYER Metal1 ;
    ANTENNADIFFAREA 2.6256 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.20115 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.098434 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 133.04996275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.995 3.155 3.935 3.155 3.935 3.01 3.835 3.01 3.835 2.69 3.935 2.69 3.935 2.07 3.995 2.07 ;
    END
  END QN
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.36 0.79 0.565 0.94 ;
    END
  END G
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.41 2.495 0.595 2.63 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 3.48 0 3.48 0 3.36 0.37 3.36 0.37 2.975 0.43 2.975 0.43 3.36 1.92 3.36 1.92 2.95 1.98 2.95 1.98 3.36 2.895 3.36 2.895 2.89 2.955 2.89 2.955 3.36 4.14 3.36 4.14 2.895 4.2 2.895 4.2 3.36 4.605 3.36 4.605 2.895 4.665 2.895 4.665 3.36 5 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5 0.06 4.67 0.06 4.67 0.545 4.61 0.545 4.61 0.06 2.54 0.06 2.54 0.49 2.48 0.49 2.48 0.06 0.385 0.06 0.385 0.495 0.325 0.495 0.325 0.06 0 0.06 0 -0.06 5 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0942 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.9074075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 33.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 0.97 1.655 1.11 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 4.495 2.755 4.405 2.755 4.405 3.155 4.345 3.155 4.345 2.07 4.405 2.07 4.405 2.695 4.495 2.695 ;
      RECT 4.3 0.4 4.36 1.365 ;
      RECT 1.445 1.485 3.71 1.545 ;
      RECT 2.155 0.7 3.31 0.76 ;
      POLYGON 3.215 2.87 3.155 2.87 3.155 1.96 2.555 1.96 2.555 1.9 3.215 1.9 ;
      POLYGON 3.065 2.82 2.645 2.82 2.645 3.035 2.585 3.035 2.585 2.875 2.37 2.875 2.37 2.815 2.585 2.815 2.585 2.76 3.005 2.76 3.005 2.125 3.065 2.125 ;
      POLYGON 2.995 0.61 2.25 0.61 2.25 0.49 2.31 0.49 2.31 0.55 2.685 0.55 2.685 0.345 2.745 0.345 2.745 0.55 2.995 0.55 ;
      POLYGON 2.995 1.23 2.745 1.23 2.745 1.305 2.685 1.305 2.685 1.09 2.745 1.09 2.745 1.17 2.995 1.17 ;
      POLYGON 2.54 1.395 2.375 1.395 2.375 1.42 2.315 1.42 2.315 1.3 2.375 1.3 2.375 1.335 2.48 1.335 2.48 1.09 2.54 1.09 ;
      POLYGON 2.29 1.2 2.08 1.2 2.08 1.305 2.02 1.305 2.02 0.355 2.08 0.355 2.08 1.14 2.29 1.14 ;
      POLYGON 2.265 2.73 2.185 2.73 2.185 3.095 2.125 3.095 2.125 2.73 2.02 2.73 2.02 2.125 2.08 2.125 2.08 2.67 2.265 2.67 ;
      POLYGON 1.875 1.335 1.21 1.335 1.21 1.275 1.815 1.275 1.815 0.355 1.875 0.355 ;
      POLYGON 1.33 2.385 0.84 2.385 0.84 3.035 0.74 3.035 0.74 3.12 0.68 3.12 0.68 2.975 0.78 2.975 0.78 2.385 0.68 2.385 0.68 2.055 0.74 2.055 0.74 2.325 1.33 2.325 ;
      POLYGON 0.985 1.1 0.69 1.1 0.69 1.385 0.63 1.385 0.63 0.495 0.53 0.495 0.53 0.35 0.59 0.35 0.59 0.435 0.69 0.435 0.69 0.7 0.92 0.7 0.92 0.76 0.69 0.76 0.69 1.04 0.985 1.04 ;
      POLYGON 0.695 2.845 0.225 2.845 0.225 3.12 0.165 3.12 0.165 2.055 0.225 2.055 0.225 2.785 0.695 2.785 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END RTLATX1

MACRO SDFF2RX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFF2RX1 0 0 ;
  SIZE 10.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.445 0.77 5.625 0.92 ;
    END
  END CK
  PIN Q2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.565075 LAYER Metal1 ;
    ANTENNADIFFAREA 9.9109 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4734 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.8679235 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 105.05703425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.14 0.96 10.09 0.96 10.09 1.11 9.96 1.11 9.96 1.05 9.995 1.05 9.995 0.54 10.07 0.54 10.07 0.6 10.075 0.6 10.075 0.76 10.14 0.76 ;
    END
  END Q2
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.565075 LAYER Metal1 ;
    ANTENNADIFFAREA 8.50985 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4734 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.8679235 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 105.05703425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.74 1.11 10.61 1.11 10.61 1.05 10.645 1.05 10.645 0.54 10.74 0.54 ;
    END
  END Q2N
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.14 0.875 7.06 0.875 7.06 0.775 7.015 0.775 7.015 0.62 7.14 0.62 ;
    END
  END D2
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.74135 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0648 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.4405865 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 108.611111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.735 1.35 7.735 1.35 7.735 1.375 7.335 1.375 7.335 1.35 6.825 1.35 6.825 1.48 6.645 1.48 6.645 1.35 3.465 1.35 3.465 1.375 3.065 1.375 3.065 1.35 0.065 1.35 0.065 1.29 3.125 1.29 3.125 1.315 3.41 1.315 3.41 1.29 7.39 1.29 7.39 1.315 7.675 1.315 7.675 1.29 10.735 1.29 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0648 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 60.83333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.735 0.41 6.57 0.41 6.57 0.7 6.835 0.7 6.835 0.865 6.775 0.865 6.775 0.76 6.51 0.76 6.51 0.41 6.145 0.41 6.145 0.895 6.06 0.895 6.06 0.41 4.74 0.41 4.74 0.895 4.655 0.895 4.655 0.41 4.29 0.41 4.29 0.76 4.025 0.76 4.025 0.865 3.965 0.865 3.965 0.7 4.23 0.7 4.23 0.41 0.065 0.41 0.065 0.35 10.735 0.35 ;
    END
  END SE
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.565075 LAYER Metal1 ;
    ANTENNADIFFAREA 8.481125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4734 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.8679235 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 105.05703425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.84 1.11 0.71 1.11 0.71 0.96 0.66 0.96 0.66 0.76 0.725 0.76 0.725 0.6 0.73 0.6 0.73 0.54 0.805 0.54 0.805 1.05 0.84 1.05 ;
    END
  END Q1
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.565075 LAYER Metal1 ;
    ANTENNADIFFAREA 8.50985 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4734 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.8679235 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 105.05703425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.19 1.11 0.06 1.11 0.06 0.54 0.155 0.54 0.155 1.05 0.19 1.05 ;
    END
  END Q1N
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.785 0.775 3.74 0.775 3.74 0.875 3.66 0.875 3.66 0.62 3.785 0.62 ;
    END
  END D1
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.39 0.625 4.565 0.77 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.8 1.77 0 1.77 0 1.65 0.3 1.65 0.3 1.54 0.42 1.54 0.42 1.65 0.955 1.65 0.955 1.54 1.075 1.54 1.075 1.65 1.53 1.65 1.53 1.54 1.65 1.54 1.65 1.65 2.445 1.65 2.445 1.54 2.565 1.54 2.565 1.65 2.795 1.65 2.795 1.54 2.915 1.54 2.915 1.65 3.675 1.65 3.675 1.54 3.795 1.54 3.795 1.65 4.465 1.65 4.465 1.54 4.585 1.54 4.585 1.65 5.33 1.65 5.33 1.54 5.45 1.54 5.45 1.65 6.215 1.65 6.215 1.54 6.335 1.54 6.335 1.65 7.005 1.65 7.005 1.54 7.125 1.54 7.125 1.65 7.885 1.65 7.885 1.54 8.005 1.54 8.005 1.65 8.235 1.65 8.235 1.54 8.355 1.54 8.355 1.65 9.15 1.65 9.15 1.54 9.27 1.54 9.27 1.65 9.725 1.65 9.725 1.54 9.845 1.54 9.845 1.65 10.38 1.65 10.38 1.54 10.5 1.54 10.5 1.65 10.8 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.8 0.06 10.5 0.06 10.5 0.17 10.38 0.17 10.38 0.06 9.895 0.06 9.895 0.17 9.775 0.17 9.775 0.06 9.27 0.06 9.27 0.17 9.15 0.17 9.15 0.06 8.255 0.06 8.255 0.17 8.135 0.17 8.135 0.06 7.15 0.06 7.15 0.17 7.03 0.17 7.03 0.06 6.335 0.06 6.335 0.17 6.215 0.17 6.215 0.06 5.45 0.06 5.45 0.17 5.325 0.17 5.325 0.06 4.585 0.06 4.585 0.17 4.465 0.17 4.465 0.06 3.77 0.06 3.77 0.17 3.65 0.17 3.65 0.06 2.665 0.06 2.665 0.17 2.545 0.17 2.545 0.06 1.65 0.06 1.65 0.17 1.53 0.17 1.53 0.06 1.025 0.06 1.025 0.17 0.905 0.17 0.905 0.06 0.42 0.06 0.42 0.17 0.3 0.17 0.3 0.06 0 0.06 0 -0.06 10.8 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 10.735 0.29 0.065 0.29 0.065 0.23 4.66 0.23 4.66 0.205 4.8 0.205 4.8 0.23 6 0.23 6 0.205 6.14 0.205 6.14 0.23 10.735 0.23 ;
      POLYGON 10.735 1.23 7.615 1.23 7.615 1.255 7.45 1.255 7.45 1.23 3.35 1.23 3.35 1.255 3.185 1.255 3.185 1.23 0.065 1.23 0.065 1.17 1.835 1.17 1.835 0.665 1.895 0.665 1.895 1.17 2.165 1.17 2.165 0.865 2.105 0.865 2.105 0.805 2.225 0.805 2.225 1.17 4.64 1.17 4.64 1.15 4.78 1.15 4.78 1.17 5.295 1.17 5.295 0.895 5.26 0.895 5.26 0.495 5.36 0.495 5.36 0.625 5.565 0.625 5.565 0.505 5.625 0.505 5.625 0.705 5.36 0.705 5.36 1.005 5.655 1.005 5.655 1.065 5.36 1.065 5.36 1.17 6.02 1.17 6.02 1.15 6.16 1.15 6.16 1.17 8.575 1.17 8.575 0.805 8.695 0.805 8.695 0.865 8.635 0.865 8.635 1.17 8.905 1.17 8.905 0.665 8.965 0.665 8.965 1.17 10.735 1.17 ;
      POLYGON 10.73 1.48 7.84 1.48 7.84 1.495 7.22 1.495 7.22 1.48 7.005 1.48 7.005 1.42 7.275 1.42 7.275 1.435 7.78 1.435 7.78 1.42 10.73 1.42 ;
      POLYGON 10.545 0.84 10.29 0.84 10.29 1.02 10.21 1.02 10.21 0.54 10.29 0.54 10.29 0.76 10.545 0.76 ;
      POLYGON 9.925 0.82 9.645 0.82 9.645 1.1 9.075 1.1 9.075 0.68 9.135 0.68 9.135 1.04 9.585 1.04 9.585 0.485 9.645 0.485 9.645 0.76 9.925 0.76 ;
      POLYGON 9.515 0.825 9.455 0.825 9.455 0.66 9.4 0.66 9.4 0.575 8.82 0.575 8.82 1.055 8.76 1.055 8.76 0.575 8.71 0.575 8.71 0.495 9.46 0.495 9.46 0.6 9.515 0.6 ;
      RECT 9.235 0.735 9.395 0.96 ;
      POLYGON 8.54 0.575 8.51 0.575 8.51 1.055 8.45 1.055 8.45 0.74 7.855 0.74 7.855 0.68 8.45 0.68 8.45 0.575 8.42 0.575 8.42 0.515 8.54 0.515 ;
      POLYGON 8.37 0.86 7.52 0.86 7.52 1.045 7.46 1.045 7.46 0.8 7.645 0.8 7.645 0.575 7.61 0.575 7.61 0.515 7.74 0.515 7.74 0.575 7.705 0.575 7.705 0.8 8.37 0.8 ;
      RECT 7.635 0.95 8.135 1.03 ;
      POLYGON 7.53 0.575 7.5 0.575 7.5 0.73 7.4 0.73 7.4 0.95 7.315 0.95 7.315 1.065 6.615 1.065 6.615 1.005 6.895 1.005 6.895 0.54 6.655 0.54 6.655 0.48 6.955 0.48 6.955 1.005 7.255 1.005 7.255 0.89 7.34 0.89 7.34 0.67 7.44 0.67 7.44 0.575 7.41 0.575 7.41 0.515 7.53 0.515 ;
      POLYGON 6.67 0.905 6.315 0.905 6.315 1.065 5.925 1.065 5.925 0.51 5.985 0.51 5.985 1.005 6.255 1.005 6.255 0.845 6.67 0.845 ;
      POLYGON 6.495 1.48 3.58 1.48 3.58 1.495 2.96 1.495 2.96 1.48 0.07 1.48 0.07 1.42 3.02 1.42 3.02 1.435 3.525 1.435 3.525 1.42 6.495 1.42 ;
      RECT 6.235 0.625 6.41 0.77 ;
      POLYGON 5.2 1.1 5.06 1.1 5.06 0.77 5.14 0.77 5.14 0.495 5.2 0.495 ;
      POLYGON 4.875 1.065 4.485 1.065 4.485 0.905 4.13 0.905 4.13 0.845 4.545 0.845 4.545 1.005 4.815 1.005 4.815 0.51 4.875 0.51 ;
      POLYGON 4.185 1.065 3.485 1.065 3.485 0.95 3.4 0.95 3.4 0.73 3.3 0.73 3.3 0.575 3.27 0.575 3.27 0.515 3.39 0.515 3.39 0.575 3.36 0.575 3.36 0.67 3.46 0.67 3.46 0.89 3.545 0.89 3.545 1.005 3.845 1.005 3.845 0.48 4.145 0.48 4.145 0.54 3.905 0.54 3.905 1.005 4.185 1.005 ;
      POLYGON 3.34 1.045 3.28 1.045 3.28 0.86 2.43 0.86 2.43 0.8 3.095 0.8 3.095 0.575 3.06 0.575 3.06 0.515 3.19 0.515 3.19 0.575 3.155 0.575 3.155 0.8 3.34 0.8 ;
      RECT 2.665 0.95 3.165 1.03 ;
      POLYGON 2.945 0.74 2.35 0.74 2.35 1.055 2.29 1.055 2.29 0.575 2.26 0.575 2.26 0.515 2.38 0.515 2.38 0.575 2.35 0.575 2.35 0.68 2.945 0.68 ;
      POLYGON 2.09 0.575 2.04 0.575 2.04 1.055 1.98 1.055 1.98 0.575 1.4 0.575 1.4 0.66 1.345 0.66 1.345 0.825 1.285 0.825 1.285 0.6 1.34 0.6 1.34 0.495 2.09 0.495 ;
      POLYGON 1.725 1.1 1.155 1.1 1.155 0.82 0.875 0.82 0.875 0.76 1.155 0.76 1.155 0.485 1.215 0.485 1.215 1.04 1.665 1.04 1.665 0.68 1.725 0.68 ;
      RECT 1.405 0.735 1.565 0.96 ;
      POLYGON 0.59 1.02 0.51 1.02 0.51 0.84 0.255 0.84 0.255 0.76 0.51 0.76 0.51 0.54 0.59 0.54 ;
  END
END SDFF2RX1

MACRO SDFF2RX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFF2RX2 0 0 ;
  SIZE 12 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.045 0.77 6.225 0.92 ;
    END
  END CK
  PIN Q2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.769075 LAYER Metal1 ;
    ANTENNADIFFAREA 10.1158 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.60435 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.2005875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.79424175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.585 0.54 10.74 1.11 ;
    END
  END Q2
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.769075 LAYER Metal1 ;
    ANTENNADIFFAREA 9.8026 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.60435 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.2005875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.79424175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.455 0.54 11.595 1.11 ;
    END
  END Q2N
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.74 0.875 7.66 0.875 7.66 0.775 7.615 0.775 7.615 0.62 7.74 0.62 ;
    END
  END D2
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.61605 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.07875 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.82285725 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 73.295238 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.28 1.35 8.335 1.35 8.335 1.375 7.935 1.375 7.935 1.35 7.44 1.35 7.44 1.48 7.25 1.48 7.25 1.35 4.065 1.35 4.065 1.375 3.665 1.375 3.665 1.35 1.72 1.35 1.72 1.29 3.725 1.29 3.725 1.315 4.01 1.315 4.01 1.29 7.99 1.29 7.99 1.315 8.275 1.315 8.275 1.29 10.28 1.29 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0648 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 51.06481475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.28 0.41 7.17 0.41 7.17 0.7 7.435 0.7 7.435 0.865 7.375 0.865 7.375 0.76 7.11 0.76 7.11 0.41 6.745 0.41 6.745 0.895 6.66 0.895 6.66 0.41 5.34 0.41 5.34 0.895 5.255 0.895 5.255 0.41 4.89 0.41 4.89 0.76 4.625 0.76 4.625 0.865 4.565 0.865 4.565 0.7 4.83 0.7 4.83 0.41 1.72 0.41 1.72 0.35 10.28 0.35 ;
    END
  END SE
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.769075 LAYER Metal1 ;
    ANTENNADIFFAREA 9.749275 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.60435 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.2005875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.79424175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.54 1.415 1.11 ;
    END
  END Q1
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.769075 LAYER Metal1 ;
    ANTENNADIFFAREA 9.8026 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.60435 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.2005875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.79424175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.405 0.54 0.545 1.11 ;
    END
  END Q1N
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.385 0.775 4.34 0.775 4.34 0.875 4.26 0.875 4.26 0.62 4.385 0.62 ;
    END
  END D1
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.99 0.625 5.165 0.77 ;
    END
  END SI
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 12 1.77 0 1.77 0 1.65 0.24 1.65 0.24 1.54 0.36 1.54 0.36 1.65 0.61 1.65 0.61 1.54 0.765 1.54 0.765 1.65 1.065 1.65 1.065 1.54 1.185 1.54 1.185 1.65 1.555 1.65 1.555 1.54 1.675 1.54 1.675 1.65 2.13 1.65 2.13 1.54 2.25 1.54 2.25 1.65 3.045 1.65 3.045 1.54 3.165 1.54 3.165 1.65 3.395 1.65 3.395 1.54 3.515 1.54 3.515 1.65 4.275 1.65 4.275 1.54 4.395 1.54 4.395 1.65 5.065 1.65 5.065 1.54 5.185 1.54 5.185 1.65 5.93 1.65 5.93 1.54 6.05 1.54 6.05 1.65 6.815 1.65 6.815 1.54 6.935 1.54 6.935 1.65 7.605 1.65 7.605 1.54 7.725 1.54 7.725 1.65 8.485 1.65 8.485 1.54 8.605 1.54 8.605 1.65 8.835 1.65 8.835 1.54 8.955 1.54 8.955 1.65 9.75 1.65 9.75 1.54 9.87 1.54 9.87 1.65 10.325 1.65 10.325 1.54 10.445 1.54 10.445 1.65 10.815 1.65 10.815 1.54 10.935 1.54 10.935 1.65 11.235 1.65 11.235 1.54 11.39 1.54 11.39 1.65 11.64 1.65 11.64 1.54 11.76 1.54 11.76 1.65 12 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 12 0.06 11.76 0.06 11.76 0.17 11.64 0.17 11.64 0.06 11.39 0.06 11.39 0.17 11.27 0.17 11.27 0.06 10.935 0.06 10.935 0.17 10.815 0.17 10.815 0.06 10.495 0.06 10.495 0.17 10.375 0.17 10.375 0.06 9.87 0.06 9.87 0.17 9.75 0.17 9.75 0.06 8.855 0.06 8.855 0.17 8.735 0.17 8.735 0.06 7.75 0.06 7.75 0.17 7.63 0.17 7.63 0.06 6.935 0.06 6.935 0.17 6.815 0.17 6.815 0.06 6.05 0.06 6.05 0.17 5.925 0.17 5.925 0.06 5.185 0.06 5.185 0.17 5.065 0.17 5.065 0.06 4.37 0.06 4.37 0.17 4.25 0.17 4.25 0.06 3.265 0.06 3.265 0.17 3.145 0.17 3.145 0.06 2.25 0.06 2.25 0.17 2.13 0.17 2.13 0.06 1.625 0.06 1.625 0.17 1.505 0.17 1.505 0.06 1.185 0.06 1.185 0.17 1.065 0.17 1.065 0.06 0.73 0.06 0.73 0.17 0.61 0.17 0.61 0.06 0.36 0.06 0.36 0.17 0.24 0.17 0.24 0.06 0 0.06 0 -0.06 12 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 11.37 0.85 11.31 0.85 11.31 0.82 11.145 0.82 11.145 1.02 11.065 1.02 11.065 0.54 11.145 0.54 11.145 0.76 11.31 0.76 11.31 0.725 11.37 0.725 ;
      POLYGON 10.525 0.82 10.245 0.82 10.245 1.1 9.675 1.1 9.675 0.68 9.735 0.68 9.735 1.04 10.185 1.04 10.185 0.485 10.245 0.485 10.245 0.76 10.525 0.76 ;
      POLYGON 10.28 0.29 1.72 0.29 1.72 0.23 5.26 0.23 5.26 0.205 5.4 0.205 5.4 0.23 6.6 0.23 6.6 0.205 6.74 0.205 6.74 0.23 10.28 0.23 ;
      POLYGON 10.28 1.23 8.215 1.23 8.215 1.255 8.05 1.255 8.05 1.23 3.95 1.23 3.95 1.255 3.785 1.255 3.785 1.23 1.72 1.23 1.72 1.17 2.435 1.17 2.435 0.665 2.495 0.665 2.495 1.17 2.765 1.17 2.765 0.865 2.705 0.865 2.705 0.805 2.825 0.805 2.825 1.17 5.24 1.17 5.24 1.15 5.38 1.15 5.38 1.17 5.895 1.17 5.895 0.895 5.86 0.895 5.86 0.495 5.96 0.495 5.96 0.625 6.165 0.625 6.165 0.505 6.225 0.505 6.225 0.705 5.96 0.705 5.96 1.005 6.255 1.005 6.255 1.065 5.96 1.065 5.96 1.17 6.62 1.17 6.62 1.15 6.76 1.15 6.76 1.17 9.175 1.17 9.175 0.805 9.295 0.805 9.295 0.865 9.235 0.865 9.235 1.17 9.505 1.17 9.505 0.665 9.565 0.665 9.565 1.17 10.28 1.17 ;
      POLYGON 10.275 1.48 8.44 1.48 8.44 1.495 7.82 1.495 7.82 1.48 7.605 1.48 7.605 1.42 7.875 1.42 7.875 1.435 8.38 1.435 8.38 1.42 10.275 1.42 ;
      POLYGON 10.115 0.825 10.055 0.825 10.055 0.66 10 0.66 10 0.575 9.42 0.575 9.42 1.055 9.36 1.055 9.36 0.575 9.31 0.575 9.31 0.495 10.06 0.495 10.06 0.6 10.115 0.6 ;
      RECT 9.835 0.735 9.995 0.96 ;
      POLYGON 9.14 0.575 9.11 0.575 9.11 1.055 9.05 1.055 9.05 0.74 8.455 0.74 8.455 0.68 9.05 0.68 9.05 0.575 9.02 0.575 9.02 0.515 9.14 0.515 ;
      POLYGON 8.97 0.86 8.12 0.86 8.12 1.045 8.06 1.045 8.06 0.8 8.245 0.8 8.245 0.575 8.21 0.575 8.21 0.515 8.34 0.515 8.34 0.575 8.305 0.575 8.305 0.8 8.97 0.8 ;
      RECT 8.235 0.95 8.735 1.03 ;
      POLYGON 8.13 0.575 8.1 0.575 8.1 0.73 8 0.73 8 0.95 7.915 0.95 7.915 1.065 7.215 1.065 7.215 1.005 7.495 1.005 7.495 0.54 7.255 0.54 7.255 0.48 7.555 0.48 7.555 1.005 7.855 1.005 7.855 0.89 7.94 0.89 7.94 0.67 8.04 0.67 8.04 0.575 8.01 0.575 8.01 0.515 8.13 0.515 ;
      POLYGON 7.27 0.905 6.915 0.905 6.915 1.065 6.525 1.065 6.525 0.51 6.585 0.51 6.585 1.005 6.855 1.005 6.855 0.845 7.27 0.845 ;
      POLYGON 7.095 1.48 4.18 1.48 4.18 1.495 3.56 1.495 3.56 1.48 1.28 1.48 1.28 1.42 3.62 1.42 3.62 1.435 4.125 1.435 4.125 1.42 7.095 1.42 ;
      RECT 6.835 0.625 7.01 0.77 ;
      POLYGON 5.8 1.1 5.66 1.1 5.66 0.77 5.74 0.77 5.74 0.495 5.8 0.495 ;
      POLYGON 5.475 1.065 5.085 1.065 5.085 0.905 4.73 0.905 4.73 0.845 5.145 0.845 5.145 1.005 5.415 1.005 5.415 0.51 5.475 0.51 ;
      POLYGON 4.785 1.065 4.085 1.065 4.085 0.95 4 0.95 4 0.73 3.9 0.73 3.9 0.575 3.87 0.575 3.87 0.515 3.99 0.515 3.99 0.575 3.96 0.575 3.96 0.67 4.06 0.67 4.06 0.89 4.145 0.89 4.145 1.005 4.445 1.005 4.445 0.48 4.745 0.48 4.745 0.54 4.505 0.54 4.505 1.005 4.785 1.005 ;
      POLYGON 3.94 1.045 3.88 1.045 3.88 0.86 3.03 0.86 3.03 0.8 3.695 0.8 3.695 0.575 3.66 0.575 3.66 0.515 3.79 0.515 3.79 0.575 3.755 0.575 3.755 0.8 3.94 0.8 ;
      RECT 3.265 0.95 3.765 1.03 ;
      POLYGON 3.545 0.74 2.95 0.74 2.95 1.055 2.89 1.055 2.89 0.575 2.86 0.575 2.86 0.515 2.98 0.515 2.98 0.575 2.95 0.575 2.95 0.68 3.545 0.68 ;
      POLYGON 2.69 0.575 2.64 0.575 2.64 1.055 2.58 1.055 2.58 0.575 2 0.575 2 0.66 1.945 0.66 1.945 0.825 1.885 0.825 1.885 0.6 1.94 0.6 1.94 0.495 2.69 0.495 ;
      POLYGON 2.325 1.1 1.755 1.1 1.755 0.82 1.475 0.82 1.475 0.76 1.755 0.76 1.755 0.485 1.815 0.485 1.815 1.04 2.265 1.04 2.265 0.68 2.325 0.68 ;
      RECT 2.005 0.735 2.165 0.96 ;
      POLYGON 0.935 1.02 0.855 1.02 0.855 0.82 0.69 0.82 0.69 0.85 0.63 0.85 0.63 0.725 0.69 0.725 0.69 0.76 0.855 0.76 0.855 0.54 0.935 0.54 ;
  END
END SDFF2RX2

MACRO SDFF4RX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFF4RX1 0 0 ;
  SIZE 20.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.844525 LAYER Metal1 ;
    ANTENNADIFFAREA 16.33035 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9468 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.5662495 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 103.35234475 LAYER Metal1 ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.8 1.77 0 1.77 0 1.65 0.3 1.65 0.3 1.54 0.42 1.54 0.42 1.65 0.955 1.65 0.955 1.54 1.075 1.54 1.075 1.65 1.53 1.65 1.53 1.54 1.65 1.54 1.65 1.65 2.445 1.65 2.445 1.54 2.565 1.54 2.565 1.65 2.795 1.65 2.795 1.54 2.915 1.54 2.915 1.65 3.675 1.65 3.675 1.54 3.795 1.54 3.795 1.65 4.465 1.65 4.465 1.54 4.585 1.54 4.585 1.65 5.415 1.65 5.415 1.54 5.535 1.54 5.535 1.65 6.205 1.65 6.205 1.54 6.325 1.54 6.325 1.65 7.085 1.65 7.085 1.54 7.205 1.54 7.205 1.65 7.435 1.65 7.435 1.54 7.555 1.54 7.555 1.65 8.35 1.65 8.35 1.54 8.47 1.54 8.47 1.65 8.925 1.65 8.925 1.54 9.045 1.54 9.045 1.65 9.58 1.65 9.58 1.54 9.7 1.54 9.7 1.65 10.35 1.65 10.35 1.54 10.47 1.54 10.47 1.65 11.215 1.65 11.215 1.54 11.335 1.54 11.335 1.65 12.005 1.65 12.005 1.54 12.125 1.54 12.125 1.65 12.885 1.65 12.885 1.54 13.005 1.54 13.005 1.65 13.235 1.65 13.235 1.54 13.355 1.54 13.355 1.65 14.15 1.65 14.15 1.54 14.27 1.54 14.27 1.65 14.725 1.65 14.725 1.54 14.845 1.54 14.845 1.65 15.38 1.65 15.38 1.54 15.5 1.54 15.5 1.65 16.215 1.65 16.215 1.54 16.335 1.54 16.335 1.65 17.005 1.65 17.005 1.54 17.125 1.54 17.125 1.65 17.885 1.65 17.885 1.54 18.005 1.54 18.005 1.65 18.235 1.65 18.235 1.54 18.355 1.54 18.355 1.65 19.15 1.65 19.15 1.54 19.27 1.54 19.27 1.65 19.725 1.65 19.725 1.54 19.845 1.54 19.845 1.65 20.38 1.65 20.38 1.54 20.5 1.54 20.5 1.65 20.8 1.65 ;
    END
  END VDD
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.175 0.77 10.355 0.92 ;
    END
  END CK
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.844525 LAYER Metal1 ;
    ANTENNADIFFAREA 13.700575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9468 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.5662495 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 103.35234475 LAYER Metal1 ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.8 0.06 20.5 0.06 20.5 0.17 20.38 0.17 20.38 0.06 19.895 0.06 19.895 0.17 19.775 0.17 19.775 0.06 19.27 0.06 19.27 0.17 19.15 0.17 19.15 0.06 18.255 0.06 18.255 0.17 18.135 0.17 18.135 0.06 17.15 0.06 17.15 0.17 17.03 0.17 17.03 0.06 16.335 0.06 16.335 0.17 16.215 0.17 16.215 0.06 15.5 0.06 15.5 0.17 15.38 0.17 15.38 0.06 14.895 0.06 14.895 0.17 14.775 0.17 14.775 0.06 14.27 0.06 14.27 0.17 14.15 0.17 14.15 0.06 13.255 0.06 13.255 0.17 13.135 0.17 13.135 0.06 12.15 0.06 12.15 0.17 12.03 0.17 12.03 0.06 11.335 0.06 11.335 0.17 11.215 0.17 11.215 0.06 10.475 0.06 10.475 0.17 10.35 0.17 10.35 0.06 9.7 0.06 9.7 0.17 9.58 0.17 9.58 0.06 9.095 0.06 9.095 0.17 8.975 0.17 8.975 0.06 8.47 0.06 8.47 0.17 8.35 0.17 8.35 0.06 7.455 0.06 7.455 0.17 7.335 0.17 7.335 0.06 6.35 0.06 6.35 0.17 6.23 0.17 6.23 0.06 5.535 0.06 5.535 0.17 5.415 0.17 5.415 0.06 4.585 0.06 4.585 0.17 4.465 0.17 4.465 0.06 3.77 0.06 3.77 0.17 3.65 0.17 3.65 0.06 2.665 0.06 2.665 0.17 2.545 0.17 2.545 0.06 1.65 0.06 1.65 0.17 1.53 0.17 1.53 0.06 1.025 0.06 1.025 0.17 0.905 0.17 0.905 0.06 0.42 0.06 0.42 0.17 0.3 0.17 0.3 0.06 0 0.06 0 -0.06 20.8 -0.06 ;
    END
  END VSS
  PIN Q2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.844525 LAYER Metal1 ;
    ANTENNADIFFAREA 16.268675 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9468 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.5662495 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 103.35234475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.34 0.96 9.29 0.96 9.29 1.11 9.16 1.11 9.16 1.05 9.195 1.05 9.195 0.54 9.27 0.54 9.27 0.6 9.275 0.6 9.275 0.76 9.34 0.76 ;
    END
  END Q2
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.844525 LAYER Metal1 ;
    ANTENNADIFFAREA 16.2974 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9468 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.5662495 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 103.35234475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.94 1.11 9.81 1.11 9.81 1.05 9.845 1.05 9.845 0.54 9.94 0.54 ;
    END
  END Q2N
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.34 0.875 6.26 0.875 6.26 0.775 6.215 0.775 6.215 0.62 6.34 0.62 ;
    END
  END D2
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.4087 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1296 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.86959875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 104.62962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.735 1.35 17.735 1.35 17.735 1.375 17.335 1.375 17.335 1.35 12.735 1.35 12.735 1.375 12.335 1.375 12.335 1.35 6.935 1.35 6.935 1.375 6.535 1.375 6.535 1.35 5.96 1.35 5.96 1.48 5.86 1.48 5.86 1.35 3.465 1.35 3.465 1.375 3.065 1.375 3.065 1.35 0.065 1.35 0.065 1.29 3.125 1.29 3.125 1.315 3.41 1.315 3.41 1.29 6.59 1.29 6.59 1.315 6.875 1.315 6.875 1.29 12.39 1.29 12.39 1.315 12.675 1.315 12.675 1.29 17.39 1.29 17.39 1.315 17.675 1.315 17.675 1.29 20.735 1.29 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1296 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 59.1435185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.735 0.41 16.57 0.41 16.57 0.7 16.835 0.7 16.835 0.865 16.775 0.865 16.775 0.76 16.51 0.76 16.51 0.41 16.145 0.41 16.145 0.895 16.06 0.895 16.06 0.41 11.57 0.41 11.57 0.7 11.835 0.7 11.835 0.865 11.775 0.865 11.775 0.76 11.51 0.76 11.51 0.41 11.145 0.41 11.145 0.895 11.06 0.895 11.06 0.41 5.77 0.41 5.77 0.7 6.035 0.7 6.035 0.865 5.975 0.865 5.975 0.76 5.71 0.76 5.71 0.41 5.345 0.41 5.345 0.895 5.26 0.895 5.26 0.41 4.74 0.41 4.74 0.895 4.655 0.895 4.655 0.41 4.29 0.41 4.29 0.76 4.025 0.76 4.025 0.865 3.965 0.865 3.965 0.7 4.23 0.7 4.23 0.41 0.065 0.41 0.065 0.35 20.735 0.35 ;
    END
  END SE
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.844525 LAYER Metal1 ;
    ANTENNADIFFAREA 16.268675 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9468 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.5662495 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 103.35234475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.84 1.11 0.71 1.11 0.71 0.96 0.66 0.96 0.66 0.76 0.725 0.76 0.725 0.6 0.73 0.6 0.73 0.54 0.805 0.54 0.805 1.05 0.84 1.05 ;
    END
  END Q1
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.844525 LAYER Metal1 ;
    ANTENNADIFFAREA 16.2974 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9468 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.5662495 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 103.35234475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.19 1.11 0.06 1.11 0.06 0.54 0.155 0.54 0.155 1.05 0.19 1.05 ;
    END
  END Q1N
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.785 0.775 3.74 0.775 3.74 0.875 3.66 0.875 3.66 0.62 3.785 0.62 ;
    END
  END D1
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.39 0.625 4.565 0.77 ;
    END
  END SI
  PIN Q4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.844525 LAYER Metal1 ;
    ANTENNADIFFAREA 18.89845 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9468 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.5662495 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 103.35234475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.14 0.96 20.09 0.96 20.09 1.11 19.96 1.11 19.96 1.05 19.995 1.05 19.995 0.54 20.07 0.54 20.07 0.6 20.075 0.6 20.075 0.76 20.14 0.76 ;
    END
  END Q4
  PIN Q4N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.844525 LAYER Metal1 ;
    ANTENNADIFFAREA 16.2974 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9468 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.5662495 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 103.35234475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.74 1.11 20.61 1.11 20.61 1.05 20.645 1.05 20.645 0.54 20.74 0.54 ;
    END
  END Q4N
  PIN D4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.14 0.875 17.06 0.875 17.06 0.775 17.015 0.775 17.015 0.62 17.14 0.62 ;
    END
  END D4
  PIN Q3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.844525 LAYER Metal1 ;
    ANTENNADIFFAREA 16.268675 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9468 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.5662495 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 103.35234475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.14 0.96 15.09 0.96 15.09 1.11 14.96 1.11 14.96 1.05 14.995 1.05 14.995 0.54 15.07 0.54 15.07 0.6 15.075 0.6 15.075 0.76 15.14 0.76 ;
    END
  END Q3
  PIN Q3N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.844525 LAYER Metal1 ;
    ANTENNADIFFAREA 16.2974 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.9468 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.5662495 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 103.35234475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.74 1.11 15.61 1.11 15.61 1.05 15.645 1.05 15.645 0.54 15.74 0.54 ;
    END
  END Q3N
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.14 0.875 12.06 0.875 12.06 0.775 12.015 0.775 12.015 0.62 12.14 0.62 ;
    END
  END D3
  OBS
    LAYER Metal1 ;
      POLYGON 20.735 0.29 0.065 0.29 0.065 0.23 4.66 0.23 4.66 0.205 4.8 0.205 4.8 0.23 5.2 0.23 5.2 0.205 5.34 0.205 5.34 0.23 11 0.23 11 0.205 11.14 0.205 11.14 0.23 16 0.23 16 0.205 16.14 0.205 16.14 0.23 20.735 0.23 ;
      POLYGON 20.735 1.23 17.615 1.23 17.615 1.255 17.45 1.255 17.45 1.23 12.615 1.23 12.615 1.255 12.45 1.255 12.45 1.23 6.815 1.23 6.815 1.255 6.65 1.255 6.65 1.23 3.35 1.23 3.35 1.255 3.185 1.255 3.185 1.23 0.065 1.23 0.065 1.17 1.835 1.17 1.835 0.665 1.895 0.665 1.895 1.17 2.165 1.17 2.165 0.865 2.105 0.865 2.105 0.805 2.225 0.805 2.225 1.17 4.64 1.17 4.64 1.15 4.78 1.15 4.78 1.17 5.22 1.17 5.22 1.15 5.36 1.15 5.36 1.17 7.775 1.17 7.775 0.805 7.895 0.805 7.895 0.865 7.835 0.865 7.835 1.17 8.105 1.17 8.105 0.665 8.165 0.665 8.165 1.17 10.44 1.17 10.44 1.065 10.145 1.065 10.145 1.005 10.44 1.005 10.44 0.705 10.175 0.705 10.175 0.505 10.235 0.505 10.235 0.625 10.44 0.625 10.44 0.495 10.54 0.495 10.54 0.895 10.505 0.895 10.505 1.17 11.02 1.17 11.02 1.15 11.16 1.15 11.16 1.17 13.575 1.17 13.575 0.805 13.695 0.805 13.695 0.865 13.635 0.865 13.635 1.17 13.905 1.17 13.905 0.665 13.965 0.665 13.965 1.17 16.02 1.17 16.02 1.15 16.16 1.15 16.16 1.17 18.575 1.17 18.575 0.805 18.695 0.805 18.695 0.865 18.635 0.865 18.635 1.17 18.905 1.17 18.905 0.665 18.965 0.665 18.965 1.17 20.735 1.17 ;
      POLYGON 20.73 1.48 17.84 1.48 17.84 1.495 17.22 1.495 17.22 1.48 17.005 1.48 17.005 1.42 17.275 1.42 17.275 1.435 17.78 1.435 17.78 1.42 20.73 1.42 ;
      POLYGON 20.545 0.84 20.29 0.84 20.29 1.02 20.21 1.02 20.21 0.54 20.29 0.54 20.29 0.76 20.545 0.76 ;
      POLYGON 19.925 0.82 19.645 0.82 19.645 1.1 19.075 1.1 19.075 0.68 19.135 0.68 19.135 1.04 19.585 1.04 19.585 0.485 19.645 0.485 19.645 0.76 19.925 0.76 ;
      POLYGON 19.515 0.825 19.455 0.825 19.455 0.66 19.4 0.66 19.4 0.575 18.82 0.575 18.82 1.055 18.76 1.055 18.76 0.575 18.71 0.575 18.71 0.495 19.46 0.495 19.46 0.6 19.515 0.6 ;
      RECT 19.235 0.735 19.395 0.96 ;
      POLYGON 18.54 0.575 18.51 0.575 18.51 1.055 18.45 1.055 18.45 0.74 17.855 0.74 17.855 0.68 18.45 0.68 18.45 0.575 18.42 0.575 18.42 0.515 18.54 0.515 ;
      POLYGON 18.37 0.86 17.52 0.86 17.52 1.045 17.46 1.045 17.46 0.8 17.645 0.8 17.645 0.575 17.61 0.575 17.61 0.515 17.74 0.515 17.74 0.575 17.705 0.575 17.705 0.8 18.37 0.8 ;
      RECT 17.635 0.95 18.135 1.03 ;
      POLYGON 17.53 0.575 17.5 0.575 17.5 0.73 17.4 0.73 17.4 0.95 17.315 0.95 17.315 1.065 16.615 1.065 16.615 1.005 16.895 1.005 16.895 0.54 16.655 0.54 16.655 0.48 16.955 0.48 16.955 1.005 17.255 1.005 17.255 0.89 17.34 0.89 17.34 0.67 17.44 0.67 17.44 0.575 17.41 0.575 17.41 0.515 17.53 0.515 ;
      POLYGON 16.67 0.905 16.315 0.905 16.315 1.065 15.925 1.065 15.925 0.51 15.985 0.51 15.985 1.005 16.255 1.005 16.255 0.845 16.67 0.845 ;
      POLYGON 16.495 1.48 12.84 1.48 12.84 1.495 12.22 1.495 12.22 1.48 12.005 1.48 12.005 1.42 12.275 1.42 12.275 1.435 12.78 1.435 12.78 1.42 16.495 1.42 ;
      RECT 16.235 0.625 16.41 0.77 ;
      POLYGON 15.545 0.84 15.29 0.84 15.29 1.02 15.21 1.02 15.21 0.54 15.29 0.54 15.29 0.76 15.545 0.76 ;
      POLYGON 14.925 0.82 14.645 0.82 14.645 1.1 14.075 1.1 14.075 0.68 14.135 0.68 14.135 1.04 14.585 1.04 14.585 0.485 14.645 0.485 14.645 0.76 14.925 0.76 ;
      POLYGON 14.515 0.825 14.455 0.825 14.455 0.66 14.4 0.66 14.4 0.575 13.82 0.575 13.82 1.055 13.76 1.055 13.76 0.575 13.71 0.575 13.71 0.495 14.46 0.495 14.46 0.6 14.515 0.6 ;
      RECT 14.235 0.735 14.395 0.96 ;
      POLYGON 13.54 0.575 13.51 0.575 13.51 1.055 13.45 1.055 13.45 0.74 12.855 0.74 12.855 0.68 13.45 0.68 13.45 0.575 13.42 0.575 13.42 0.515 13.54 0.515 ;
      POLYGON 13.37 0.86 12.52 0.86 12.52 1.045 12.46 1.045 12.46 0.8 12.645 0.8 12.645 0.575 12.61 0.575 12.61 0.515 12.74 0.515 12.74 0.575 12.705 0.575 12.705 0.8 13.37 0.8 ;
      RECT 12.635 0.95 13.135 1.03 ;
      POLYGON 12.53 0.575 12.5 0.575 12.5 0.73 12.4 0.73 12.4 0.95 12.315 0.95 12.315 1.065 11.615 1.065 11.615 1.005 11.895 1.005 11.895 0.54 11.655 0.54 11.655 0.48 11.955 0.48 11.955 1.005 12.255 1.005 12.255 0.89 12.34 0.89 12.34 0.67 12.44 0.67 12.44 0.575 12.41 0.575 12.41 0.515 12.53 0.515 ;
      POLYGON 11.67 0.905 11.315 0.905 11.315 1.065 10.925 1.065 10.925 0.51 10.985 0.51 10.985 1.005 11.255 1.005 11.255 0.845 11.67 0.845 ;
      POLYGON 11.495 1.48 7.04 1.48 7.04 1.495 6.42 1.495 6.42 1.48 6.205 1.48 6.205 1.42 6.475 1.42 6.475 1.435 6.98 1.435 6.98 1.42 11.495 1.42 ;
      RECT 11.235 0.625 11.41 0.77 ;
      POLYGON 10.74 1.1 10.6 1.1 10.6 0.495 10.66 0.495 10.66 0.77 10.74 0.77 ;
      POLYGON 9.745 0.84 9.49 0.84 9.49 1.02 9.41 1.02 9.41 0.54 9.49 0.54 9.49 0.76 9.745 0.76 ;
      POLYGON 9.125 0.82 8.845 0.82 8.845 1.1 8.275 1.1 8.275 0.68 8.335 0.68 8.335 1.04 8.785 1.04 8.785 0.485 8.845 0.485 8.845 0.76 9.125 0.76 ;
      POLYGON 8.715 0.825 8.655 0.825 8.655 0.66 8.6 0.66 8.6 0.575 8.02 0.575 8.02 1.055 7.96 1.055 7.96 0.575 7.91 0.575 7.91 0.495 8.66 0.495 8.66 0.6 8.715 0.6 ;
      RECT 8.435 0.735 8.595 0.96 ;
      POLYGON 7.74 0.575 7.71 0.575 7.71 1.055 7.65 1.055 7.65 0.74 7.055 0.74 7.055 0.68 7.65 0.68 7.65 0.575 7.62 0.575 7.62 0.515 7.74 0.515 ;
      POLYGON 7.57 0.86 6.72 0.86 6.72 1.045 6.66 1.045 6.66 0.8 6.845 0.8 6.845 0.575 6.81 0.575 6.81 0.515 6.94 0.515 6.94 0.575 6.905 0.575 6.905 0.8 7.57 0.8 ;
      RECT 6.835 0.95 7.335 1.03 ;
      POLYGON 6.73 0.575 6.7 0.575 6.7 0.73 6.6 0.73 6.6 0.95 6.515 0.95 6.515 1.065 5.815 1.065 5.815 1.005 6.095 1.005 6.095 0.54 5.855 0.54 5.855 0.48 6.155 0.48 6.155 1.005 6.455 1.005 6.455 0.89 6.54 0.89 6.54 0.67 6.64 0.67 6.64 0.575 6.61 0.575 6.61 0.515 6.73 0.515 ;
      POLYGON 5.87 0.905 5.515 0.905 5.515 1.065 5.125 1.065 5.125 0.51 5.185 0.51 5.185 1.005 5.455 1.005 5.455 0.845 5.87 0.845 ;
      POLYGON 5.695 1.48 3.58 1.48 3.58 1.495 2.96 1.495 2.96 1.48 0.07 1.48 0.07 1.42 3.02 1.42 3.02 1.435 3.525 1.435 3.525 1.42 5.695 1.42 ;
      RECT 5.435 0.625 5.61 0.77 ;
      POLYGON 4.875 1.065 4.485 1.065 4.485 0.905 4.13 0.905 4.13 0.845 4.545 0.845 4.545 1.005 4.815 1.005 4.815 0.51 4.875 0.51 ;
      POLYGON 4.185 1.065 3.485 1.065 3.485 0.95 3.4 0.95 3.4 0.73 3.3 0.73 3.3 0.575 3.27 0.575 3.27 0.515 3.39 0.515 3.39 0.575 3.36 0.575 3.36 0.67 3.46 0.67 3.46 0.89 3.545 0.89 3.545 1.005 3.845 1.005 3.845 0.48 4.145 0.48 4.145 0.54 3.905 0.54 3.905 1.005 4.185 1.005 ;
      POLYGON 3.34 1.045 3.28 1.045 3.28 0.86 2.43 0.86 2.43 0.8 3.095 0.8 3.095 0.575 3.06 0.575 3.06 0.515 3.19 0.515 3.19 0.575 3.155 0.575 3.155 0.8 3.34 0.8 ;
      RECT 2.665 0.95 3.165 1.03 ;
      POLYGON 2.945 0.74 2.35 0.74 2.35 1.055 2.29 1.055 2.29 0.575 2.26 0.575 2.26 0.515 2.38 0.515 2.38 0.575 2.35 0.575 2.35 0.68 2.945 0.68 ;
      POLYGON 2.09 0.575 2.04 0.575 2.04 1.055 1.98 1.055 1.98 0.575 1.4 0.575 1.4 0.66 1.345 0.66 1.345 0.825 1.285 0.825 1.285 0.6 1.34 0.6 1.34 0.495 2.09 0.495 ;
      POLYGON 1.725 1.1 1.155 1.1 1.155 0.82 0.875 0.82 0.875 0.76 1.155 0.76 1.155 0.485 1.215 0.485 1.215 1.04 1.665 1.04 1.665 0.68 1.725 0.68 ;
      RECT 1.405 0.735 1.565 0.96 ;
      POLYGON 0.59 1.02 0.51 1.02 0.51 0.84 0.255 0.84 0.255 0.76 0.51 0.76 0.51 0.54 0.59 0.54 ;
  END
END SDFF4RX1

MACRO SDFF4RX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFF4RX2 0 0 ;
  SIZE 23.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.750825 LAYER Metal1 ;
    ANTENNADIFFAREA 18.74845 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.2087 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.376541 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 83.581534 LAYER Metal1 ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.2 1.77 0 1.77 0 1.65 0.24 1.65 0.24 1.54 0.36 1.54 0.36 1.65 0.61 1.65 0.61 1.54 0.765 1.54 0.765 1.65 1.065 1.65 1.065 1.54 1.185 1.54 1.185 1.65 1.555 1.65 1.555 1.54 1.675 1.54 1.675 1.65 2.13 1.65 2.13 1.54 2.25 1.54 2.25 1.65 3.045 1.65 3.045 1.54 3.165 1.54 3.165 1.65 3.395 1.65 3.395 1.54 3.515 1.54 3.515 1.65 4.275 1.65 4.275 1.54 4.395 1.54 4.395 1.65 5.065 1.65 5.065 1.54 5.185 1.54 5.185 1.65 6.015 1.65 6.015 1.54 6.135 1.54 6.135 1.65 6.805 1.65 6.805 1.54 6.925 1.54 6.925 1.65 7.685 1.65 7.685 1.54 7.805 1.54 7.805 1.65 8.035 1.65 8.035 1.54 8.155 1.54 8.155 1.65 8.95 1.65 8.95 1.54 9.07 1.54 9.07 1.65 9.525 1.65 9.525 1.54 9.645 1.54 9.645 1.65 10.015 1.65 10.015 1.54 10.135 1.54 10.135 1.65 10.435 1.65 10.435 1.54 10.59 1.54 10.59 1.65 10.84 1.65 10.84 1.54 10.96 1.54 10.96 1.65 11.55 1.65 11.55 1.54 11.67 1.54 11.67 1.65 12.415 1.65 12.415 1.54 12.535 1.54 12.535 1.65 13.205 1.65 13.205 1.54 13.325 1.54 13.325 1.65 14.085 1.65 14.085 1.54 14.205 1.54 14.205 1.65 14.435 1.65 14.435 1.54 14.555 1.54 14.555 1.65 15.35 1.65 15.35 1.54 15.47 1.54 15.47 1.65 15.925 1.65 15.925 1.54 16.045 1.54 16.045 1.65 16.415 1.65 16.415 1.54 16.535 1.54 16.535 1.65 16.835 1.65 16.835 1.54 16.99 1.54 16.99 1.65 17.24 1.65 17.24 1.54 17.36 1.54 17.36 1.65 18.015 1.65 18.015 1.54 18.135 1.54 18.135 1.65 18.805 1.65 18.805 1.54 18.925 1.54 18.925 1.65 19.685 1.65 19.685 1.54 19.805 1.54 19.805 1.65 20.035 1.65 20.035 1.54 20.155 1.54 20.155 1.65 20.95 1.65 20.95 1.54 21.07 1.54 21.07 1.65 21.525 1.65 21.525 1.54 21.645 1.54 21.645 1.65 22.015 1.65 22.015 1.54 22.135 1.54 22.135 1.65 22.435 1.65 22.435 1.54 22.59 1.54 22.59 1.65 22.84 1.65 22.84 1.54 22.96 1.54 22.96 1.65 23.2 1.65 ;
    END
  END VDD
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.375 0.77 11.555 0.92 ;
    END
  END CK
  PIN VSS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.750825 LAYER Metal1 ;
    ANTENNADIFFAREA 15.830675 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.2087 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.376541 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 83.581534 LAYER Metal1 ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.2 0.06 22.96 0.06 22.96 0.17 22.84 0.17 22.84 0.06 22.59 0.06 22.59 0.17 22.47 0.17 22.47 0.06 22.135 0.06 22.135 0.17 22.015 0.17 22.015 0.06 21.695 0.06 21.695 0.17 21.575 0.17 21.575 0.06 21.07 0.06 21.07 0.17 20.95 0.17 20.95 0.06 20.055 0.06 20.055 0.17 19.935 0.17 19.935 0.06 18.95 0.06 18.95 0.17 18.83 0.17 18.83 0.06 18.135 0.06 18.135 0.17 18.015 0.17 18.015 0.06 17.36 0.06 17.36 0.17 17.24 0.17 17.24 0.06 16.99 0.06 16.99 0.17 16.87 0.17 16.87 0.06 16.535 0.06 16.535 0.17 16.415 0.17 16.415 0.06 16.095 0.06 16.095 0.17 15.975 0.17 15.975 0.06 15.47 0.06 15.47 0.17 15.35 0.17 15.35 0.06 14.455 0.06 14.455 0.17 14.335 0.17 14.335 0.06 13.35 0.06 13.35 0.17 13.23 0.17 13.23 0.06 12.535 0.06 12.535 0.17 12.415 0.17 12.415 0.06 11.675 0.06 11.675 0.17 11.55 0.17 11.55 0.06 10.96 0.06 10.96 0.17 10.84 0.17 10.84 0.06 10.59 0.06 10.59 0.17 10.47 0.17 10.47 0.06 10.135 0.06 10.135 0.17 10.015 0.17 10.015 0.06 9.695 0.06 9.695 0.17 9.575 0.17 9.575 0.06 9.07 0.06 9.07 0.17 8.95 0.17 8.95 0.06 8.055 0.06 8.055 0.17 7.935 0.17 7.935 0.06 6.95 0.06 6.95 0.17 6.83 0.17 6.83 0.06 6.135 0.06 6.135 0.17 6.015 0.17 6.015 0.06 5.185 0.06 5.185 0.17 5.065 0.17 5.065 0.06 4.37 0.06 4.37 0.17 4.25 0.17 4.25 0.06 3.265 0.06 3.265 0.17 3.145 0.17 3.145 0.06 2.25 0.06 2.25 0.17 2.13 0.17 2.13 0.06 1.625 0.06 1.625 0.17 1.505 0.17 1.505 0.06 1.185 0.06 1.185 0.17 1.065 0.17 1.065 0.06 0.73 0.06 0.73 0.17 0.61 0.17 0.61 0.06 0.36 0.06 0.36 0.17 0.24 0.17 0.24 0.06 0 0.06 0 -0.06 23.2 -0.06 ;
    END
  END VSS
  PIN Q2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.750825 LAYER Metal1 ;
    ANTENNADIFFAREA 19.1124 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.2087 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.376541 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 83.581534 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.785 0.54 9.94 1.11 ;
    END
  END Q2
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.750825 LAYER Metal1 ;
    ANTENNADIFFAREA 18.7992 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.2087 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.376541 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 83.581534 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.655 0.54 10.795 1.11 ;
    END
  END Q2N
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.94 0.875 6.86 0.875 6.86 0.775 6.815 0.775 6.815 0.62 6.94 0.62 ;
    END
  END D2
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3579 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1575 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.62158725 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 82.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 21.48 1.35 19.535 1.35 19.535 1.375 19.135 1.375 19.135 1.35 13.935 1.35 13.935 1.375 13.535 1.375 13.535 1.35 7.535 1.35 7.535 1.375 7.135 1.375 7.135 1.35 4.065 1.35 4.065 1.375 3.665 1.375 3.665 1.35 1.72 1.35 1.72 1.29 3.725 1.29 3.725 1.315 4.01 1.315 4.01 1.29 7.19 1.29 7.19 1.315 7.475 1.315 7.475 1.29 11.05 1.29 11.05 1.15 11.17 1.15 11.17 1.29 13.59 1.29 13.59 1.315 13.875 1.315 13.875 1.29 19.19 1.29 19.19 1.315 19.475 1.315 19.475 1.29 21.48 1.29 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1296 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 57.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 21.48 0.41 18.37 0.41 18.37 0.7 18.635 0.7 18.635 0.865 18.575 0.865 18.575 0.76 18.31 0.76 18.31 0.41 17.945 0.41 17.945 0.895 17.86 0.895 17.86 0.41 12.77 0.41 12.77 0.7 13.035 0.7 13.035 0.865 12.975 0.865 12.975 0.76 12.71 0.76 12.71 0.41 12.345 0.41 12.345 0.895 12.26 0.895 12.26 0.41 6.37 0.41 6.37 0.7 6.635 0.7 6.635 0.865 6.575 0.865 6.575 0.76 6.31 0.76 6.31 0.41 5.945 0.41 5.945 0.895 5.86 0.895 5.86 0.41 5.34 0.41 5.34 0.895 5.255 0.895 5.255 0.41 4.89 0.41 4.89 0.76 4.625 0.76 4.625 0.865 4.565 0.865 4.565 0.7 4.83 0.7 4.83 0.41 1.72 0.41 1.72 0.35 21.48 0.35 ;
    END
  END SE
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.750825 LAYER Metal1 ;
    ANTENNADIFFAREA 18.745875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.2087 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.376541 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 83.581534 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.54 1.415 1.11 ;
    END
  END Q1
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.750825 LAYER Metal1 ;
    ANTENNADIFFAREA 18.7992 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.2087 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.376541 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 83.581534 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.405 0.54 0.545 1.11 ;
    END
  END Q1N
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.385 0.775 4.34 0.775 4.34 0.875 4.26 0.875 4.26 0.62 4.385 0.62 ;
    END
  END D1
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.99 0.625 5.165 0.77 ;
    END
  END SI
  PIN Q4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.750825 LAYER Metal1 ;
    ANTENNADIFFAREA 19.1124 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.2087 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.376541 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 83.581534 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 21.785 0.54 21.94 1.11 ;
    END
  END Q4
  PIN Q4N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.750825 LAYER Metal1 ;
    ANTENNADIFFAREA 18.7992 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.2087 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.376541 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 83.581534 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 22.655 0.54 22.795 1.11 ;
    END
  END Q4N
  PIN D4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.94 0.875 18.86 0.875 18.86 0.775 18.815 0.775 18.815 0.62 18.94 0.62 ;
    END
  END D4
  PIN Q3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.750825 LAYER Metal1 ;
    ANTENNADIFFAREA 19.1124 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.2087 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.376541 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 83.581534 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 16.185 0.54 16.34 1.11 ;
    END
  END Q3
  PIN Q3N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.750825 LAYER Metal1 ;
    ANTENNADIFFAREA 18.7992 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.2087 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.376541 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 83.581534 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 17.055 0.54 17.195 1.11 ;
    END
  END Q3N
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.34 0.875 13.26 0.875 13.26 0.775 13.215 0.775 13.215 0.62 13.34 0.62 ;
    END
  END D3
  OBS
    LAYER Metal1 ;
      POLYGON 22.57 0.85 22.51 0.85 22.51 0.82 22.345 0.82 22.345 1.02 22.265 1.02 22.265 0.54 22.345 0.54 22.345 0.76 22.51 0.76 22.51 0.725 22.57 0.725 ;
      POLYGON 21.725 0.82 21.445 0.82 21.445 1.1 20.875 1.1 20.875 0.68 20.935 0.68 20.935 1.04 21.385 1.04 21.385 0.485 21.445 0.485 21.445 0.76 21.725 0.76 ;
      POLYGON 21.48 0.29 1.72 0.29 1.72 0.23 5.26 0.23 5.26 0.205 5.4 0.205 5.4 0.23 5.8 0.23 5.8 0.205 5.94 0.205 5.94 0.23 12.2 0.23 12.2 0.205 12.34 0.205 12.34 0.23 17.8 0.23 17.8 0.205 17.94 0.205 17.94 0.23 21.48 0.23 ;
      POLYGON 21.48 1.23 19.415 1.23 19.415 1.255 19.25 1.255 19.25 1.23 13.815 1.23 13.815 1.255 13.65 1.255 13.65 1.23 11.64 1.23 11.64 1.065 10.945 1.065 10.945 1.23 7.415 1.23 7.415 1.255 7.25 1.255 7.25 1.23 3.95 1.23 3.95 1.255 3.785 1.255 3.785 1.23 1.72 1.23 1.72 1.17 2.435 1.17 2.435 0.665 2.495 0.665 2.495 1.17 2.765 1.17 2.765 0.865 2.705 0.865 2.705 0.805 2.825 0.805 2.825 1.17 5.24 1.17 5.24 1.15 5.38 1.15 5.38 1.17 5.82 1.17 5.82 1.15 5.96 1.15 5.96 1.17 8.375 1.17 8.375 0.805 8.495 0.805 8.495 0.865 8.435 0.865 8.435 1.17 8.705 1.17 8.705 0.665 8.765 0.665 8.765 1.17 10.885 1.17 10.885 1.005 11.64 1.005 11.64 0.705 11.375 0.705 11.375 0.505 11.435 0.505 11.435 0.625 11.64 0.625 11.64 0.495 11.74 0.495 11.74 0.895 11.705 0.895 11.705 1.17 12.22 1.17 12.22 1.15 12.36 1.15 12.36 1.17 14.775 1.17 14.775 0.805 14.895 0.805 14.895 0.865 14.835 0.865 14.835 1.17 15.105 1.17 15.105 0.665 15.165 0.665 15.165 1.17 17.82 1.17 17.82 1.15 17.96 1.15 17.96 1.17 20.375 1.17 20.375 0.805 20.495 0.805 20.495 0.865 20.435 0.865 20.435 1.17 20.705 1.17 20.705 0.665 20.765 0.665 20.765 1.17 21.48 1.17 ;
      POLYGON 21.475 1.48 19.64 1.48 19.64 1.495 19.02 1.495 19.02 1.48 18.805 1.48 18.805 1.42 19.075 1.42 19.075 1.435 19.58 1.435 19.58 1.42 21.475 1.42 ;
      POLYGON 21.315 0.825 21.255 0.825 21.255 0.66 21.2 0.66 21.2 0.575 20.62 0.575 20.62 1.055 20.56 1.055 20.56 0.575 20.51 0.575 20.51 0.495 21.26 0.495 21.26 0.6 21.315 0.6 ;
      RECT 21.035 0.735 21.195 0.96 ;
      POLYGON 20.34 0.575 20.31 0.575 20.31 1.055 20.25 1.055 20.25 0.74 19.655 0.74 19.655 0.68 20.25 0.68 20.25 0.575 20.22 0.575 20.22 0.515 20.34 0.515 ;
      POLYGON 20.17 0.86 19.32 0.86 19.32 1.045 19.26 1.045 19.26 0.8 19.445 0.8 19.445 0.575 19.41 0.575 19.41 0.515 19.54 0.515 19.54 0.575 19.505 0.575 19.505 0.8 20.17 0.8 ;
      RECT 19.435 0.95 19.935 1.03 ;
      POLYGON 19.33 0.575 19.3 0.575 19.3 0.73 19.2 0.73 19.2 0.95 19.115 0.95 19.115 1.065 18.415 1.065 18.415 1.005 18.695 1.005 18.695 0.54 18.455 0.54 18.455 0.48 18.755 0.48 18.755 1.005 19.055 1.005 19.055 0.89 19.14 0.89 19.14 0.67 19.24 0.67 19.24 0.575 19.21 0.575 19.21 0.515 19.33 0.515 ;
      POLYGON 18.47 0.905 18.115 0.905 18.115 1.065 17.725 1.065 17.725 0.51 17.785 0.51 17.785 1.005 18.055 1.005 18.055 0.845 18.47 0.845 ;
      POLYGON 18.295 1.48 14.04 1.48 14.04 1.495 13.42 1.495 13.42 1.48 13.205 1.48 13.205 1.42 13.475 1.42 13.475 1.435 13.98 1.435 13.98 1.42 18.295 1.42 ;
      RECT 18.035 0.625 18.21 0.77 ;
      POLYGON 16.97 0.85 16.91 0.85 16.91 0.82 16.745 0.82 16.745 1.02 16.665 1.02 16.665 0.54 16.745 0.54 16.745 0.76 16.91 0.76 16.91 0.725 16.97 0.725 ;
      POLYGON 16.125 0.82 15.845 0.82 15.845 1.1 15.275 1.1 15.275 0.68 15.335 0.68 15.335 1.04 15.785 1.04 15.785 0.485 15.845 0.485 15.845 0.76 16.125 0.76 ;
      POLYGON 15.715 0.825 15.655 0.825 15.655 0.66 15.6 0.66 15.6 0.575 15.02 0.575 15.02 1.055 14.96 1.055 14.96 0.575 14.91 0.575 14.91 0.495 15.66 0.495 15.66 0.6 15.715 0.6 ;
      RECT 15.435 0.735 15.595 0.96 ;
      POLYGON 14.74 0.575 14.71 0.575 14.71 1.055 14.65 1.055 14.65 0.74 14.055 0.74 14.055 0.68 14.65 0.68 14.65 0.575 14.62 0.575 14.62 0.515 14.74 0.515 ;
      POLYGON 14.57 0.86 13.72 0.86 13.72 1.045 13.66 1.045 13.66 0.8 13.845 0.8 13.845 0.575 13.81 0.575 13.81 0.515 13.94 0.515 13.94 0.575 13.905 0.575 13.905 0.8 14.57 0.8 ;
      RECT 13.835 0.95 14.335 1.03 ;
      POLYGON 13.73 0.575 13.7 0.575 13.7 0.73 13.6 0.73 13.6 0.95 13.515 0.95 13.515 1.065 12.815 1.065 12.815 1.005 13.095 1.005 13.095 0.54 12.855 0.54 12.855 0.48 13.155 0.48 13.155 1.005 13.455 1.005 13.455 0.89 13.54 0.89 13.54 0.67 13.64 0.67 13.64 0.575 13.61 0.575 13.61 0.515 13.73 0.515 ;
      POLYGON 12.87 0.905 12.515 0.905 12.515 1.065 12.125 1.065 12.125 0.51 12.185 0.51 12.185 1.005 12.455 1.005 12.455 0.845 12.87 0.845 ;
      POLYGON 12.695 1.48 7.64 1.48 7.64 1.495 7.02 1.495 7.02 1.48 6.805 1.48 6.805 1.42 7.075 1.42 7.075 1.435 7.58 1.435 7.58 1.42 12.695 1.42 ;
      RECT 12.435 0.625 12.61 0.77 ;
      POLYGON 11.94 1.1 11.8 1.1 11.8 0.495 11.86 0.495 11.86 0.77 11.94 0.77 ;
      POLYGON 10.57 0.85 10.51 0.85 10.51 0.82 10.345 0.82 10.345 1.02 10.265 1.02 10.265 0.54 10.345 0.54 10.345 0.76 10.51 0.76 10.51 0.725 10.57 0.725 ;
      POLYGON 9.725 0.82 9.445 0.82 9.445 1.1 8.875 1.1 8.875 0.68 8.935 0.68 8.935 1.04 9.385 1.04 9.385 0.485 9.445 0.485 9.445 0.76 9.725 0.76 ;
      POLYGON 9.315 0.825 9.255 0.825 9.255 0.66 9.2 0.66 9.2 0.575 8.62 0.575 8.62 1.055 8.56 1.055 8.56 0.575 8.51 0.575 8.51 0.495 9.26 0.495 9.26 0.6 9.315 0.6 ;
      RECT 9.035 0.735 9.195 0.96 ;
      POLYGON 8.34 0.575 8.31 0.575 8.31 1.055 8.25 1.055 8.25 0.74 7.655 0.74 7.655 0.68 8.25 0.68 8.25 0.575 8.22 0.575 8.22 0.515 8.34 0.515 ;
      POLYGON 8.17 0.86 7.32 0.86 7.32 1.045 7.26 1.045 7.26 0.8 7.445 0.8 7.445 0.575 7.41 0.575 7.41 0.515 7.54 0.515 7.54 0.575 7.505 0.575 7.505 0.8 8.17 0.8 ;
      RECT 7.435 0.95 7.935 1.03 ;
      POLYGON 7.33 0.575 7.3 0.575 7.3 0.73 7.2 0.73 7.2 0.95 7.115 0.95 7.115 1.065 6.415 1.065 6.415 1.005 6.695 1.005 6.695 0.54 6.455 0.54 6.455 0.48 6.755 0.48 6.755 1.005 7.055 1.005 7.055 0.89 7.14 0.89 7.14 0.67 7.24 0.67 7.24 0.575 7.21 0.575 7.21 0.515 7.33 0.515 ;
      POLYGON 6.47 0.905 6.115 0.905 6.115 1.065 5.725 1.065 5.725 0.51 5.785 0.51 5.785 1.005 6.055 1.005 6.055 0.845 6.47 0.845 ;
      POLYGON 6.295 1.48 4.18 1.48 4.18 1.495 3.56 1.495 3.56 1.48 1.275 1.48 1.275 1.42 3.62 1.42 3.62 1.435 4.125 1.435 4.125 1.42 6.295 1.42 ;
      RECT 6.035 0.625 6.21 0.77 ;
      POLYGON 5.475 1.065 5.085 1.065 5.085 0.905 4.73 0.905 4.73 0.845 5.145 0.845 5.145 1.005 5.415 1.005 5.415 0.51 5.475 0.51 ;
      POLYGON 4.785 1.065 4.085 1.065 4.085 0.95 4 0.95 4 0.73 3.9 0.73 3.9 0.575 3.87 0.575 3.87 0.515 3.99 0.515 3.99 0.575 3.96 0.575 3.96 0.67 4.06 0.67 4.06 0.89 4.145 0.89 4.145 1.005 4.445 1.005 4.445 0.48 4.745 0.48 4.745 0.54 4.505 0.54 4.505 1.005 4.785 1.005 ;
      POLYGON 3.94 1.045 3.88 1.045 3.88 0.86 3.03 0.86 3.03 0.8 3.695 0.8 3.695 0.575 3.66 0.575 3.66 0.515 3.79 0.515 3.79 0.575 3.755 0.575 3.755 0.8 3.94 0.8 ;
      RECT 3.265 0.95 3.765 1.03 ;
      POLYGON 3.545 0.74 2.95 0.74 2.95 1.055 2.89 1.055 2.89 0.575 2.86 0.575 2.86 0.515 2.98 0.515 2.98 0.575 2.95 0.575 2.95 0.68 3.545 0.68 ;
      POLYGON 2.69 0.575 2.64 0.575 2.64 1.055 2.58 1.055 2.58 0.575 2 0.575 2 0.66 1.945 0.66 1.945 0.825 1.885 0.825 1.885 0.6 1.94 0.6 1.94 0.495 2.69 0.495 ;
      POLYGON 2.325 1.1 1.755 1.1 1.755 0.82 1.475 0.82 1.475 0.76 1.755 0.76 1.755 0.485 1.815 0.485 1.815 1.04 2.265 1.04 2.265 0.68 2.325 0.68 ;
      RECT 2.005 0.735 2.165 0.96 ;
      POLYGON 0.935 1.02 0.855 1.02 0.855 0.82 0.69 0.82 0.69 0.85 0.63 0.85 0.63 0.725 0.69 0.725 0.69 0.76 0.855 0.76 0.855 0.54 0.935 0.54 ;
  END
END SDFF4RX2

MACRO SDFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFHQX1 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.616225 LAYER Metal1 ;
    ANTENNADIFFAREA 3.24895 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2601 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.05853525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 79.25605525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.2 1.475 0.14 1.475 0.14 0.73 0.06 0.73 0.06 0.6 0.14 0.6 0.14 0.54 0.2 0.54 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.88778875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.77 0.745 4.71 0.745 4.71 0.705 3.995 0.705 3.995 0.945 3.935 0.945 3.935 0.645 4.635 0.645 4.635 0.625 4.77 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.61 0.895 4.565 0.895 4.565 1.04 4.265 1.04 4.265 0.805 4.61 0.805 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.675 0.91 3.595 0.91 3.595 0.73 3.46 0.73 3.46 0.545 3.54 0.545 3.54 0.65 3.675 0.65 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.565 1.035 0.54 1.035 0.54 1.255 0.46 1.255 0.46 0.79 0.485 0.79 0.485 0.78 0.565 0.78 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 1.77 0 1.77 0 1.65 0.345 1.65 0.345 1.355 0.405 1.355 0.405 1.65 1.11 1.65 1.11 1.29 1.23 1.29 1.23 1.35 1.17 1.35 1.17 1.65 2.365 1.65 2.365 1.365 2.485 1.365 2.485 1.425 2.425 1.425 2.425 1.65 3.615 1.65 3.615 1.17 3.675 1.17 3.675 1.65 4.425 1.65 4.425 1.315 4.485 1.315 4.485 1.65 5 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 0.06 4.54 0.06 4.54 0.525 4.48 0.525 4.48 0.06 3.675 0.06 3.675 0.415 3.615 0.415 3.615 0.06 2.425 0.06 2.425 0.19 2.485 0.19 2.485 0.25 2.365 0.25 2.365 0.06 1.225 0.06 1.225 0.49 1.165 0.49 1.165 0.06 0.405 0.06 0.405 0.52 0.345 0.52 0.345 0.06 0 0.06 0 -0.06 5 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.93 1.2 4.845 1.2 4.845 1.26 4.785 1.26 4.785 1.2 4.105 1.2 4.105 0.885 4.165 0.885 4.165 1.14 4.87 1.14 4.87 0.43 4.93 0.43 ;
      POLYGON 4.23 0.545 3.835 0.545 3.835 1.045 4.005 1.045 4.005 1.435 3.945 1.435 3.945 1.105 3.775 1.105 3.775 1.07 3.21 1.07 3.21 1.13 3.15 1.13 3.15 1.01 3.21 1.01 3.21 0.545 3.15 0.545 3.15 0.485 3.27 0.485 3.27 1.01 3.775 1.01 3.775 0.485 4.17 0.485 4.17 0.425 4.23 0.425 ;
      POLYGON 3.47 1.23 3.37 1.23 3.37 1.29 2.99 1.29 2.99 0.355 2.67 0.355 2.67 0.615 2.73 0.615 2.73 0.735 2.67 0.735 2.67 0.675 2.61 0.675 2.61 0.41 2.205 0.41 2.205 0.385 1.885 0.385 1.885 0.66 1.87 0.66 1.87 0.81 1.585 0.81 1.585 0.87 1.525 0.87 1.525 0.75 1.81 0.75 1.81 0.615 1.825 0.615 1.825 0.325 2.265 0.325 2.265 0.35 2.61 0.35 2.61 0.295 3.44 0.295 3.44 0.415 3.38 0.415 3.38 0.355 3.05 0.355 3.05 1.23 3.31 1.23 3.31 1.17 3.47 1.17 ;
      POLYGON 2.89 1.205 2.83 1.205 2.83 1.005 2.29 1.005 2.29 0.755 2.35 0.755 2.35 0.945 2.83 0.945 2.83 0.515 2.77 0.515 2.77 0.455 2.89 0.455 ;
      POLYGON 2.78 1.365 2.66 1.365 2.66 1.265 1.43 1.265 1.43 1.19 0.725 1.19 0.725 1.38 0.665 1.38 0.665 0.54 0.725 0.54 0.725 1.13 1.49 1.13 1.49 1.205 1.97 1.205 1.97 0.765 2.03 0.765 2.03 1.205 2.72 1.205 2.72 1.305 2.78 1.305 ;
      POLYGON 2.51 0.845 2.45 0.845 2.45 0.655 2.19 0.655 2.19 1.105 2.13 1.105 2.13 0.57 1.985 0.57 1.985 0.485 2.105 0.485 2.105 0.51 2.19 0.51 2.19 0.595 2.51 0.595 ;
      POLYGON 1.725 0.545 1.425 0.545 1.425 0.97 1.65 0.97 1.65 1.105 1.59 1.105 1.59 1.03 1.045 1.03 1.045 0.87 1.035 0.87 1.035 0.75 1.105 0.75 1.105 0.97 1.365 0.97 1.365 0.485 1.725 0.485 ;
      POLYGON 1.265 0.865 1.205 0.865 1.205 0.65 0.885 0.65 0.885 0.97 0.945 0.97 0.945 1.03 0.825 1.03 0.825 0.44 0.565 0.44 0.565 0.68 0.36 0.68 0.36 0.82 0.3 0.82 0.3 0.62 0.505 0.62 0.505 0.38 1.02 0.38 1.02 0.59 1.265 0.59 ;
  END
END SDFFHQX1

MACRO SDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFHQX2 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.763325 LAYER Metal1 ;
    ANTENNADIFFAREA 3.4928 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.28935 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.55011225 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 74.88335925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.36 1.335 0.3 1.335 0.3 0.92 0.26 0.92 0.26 0.79 0.3 0.79 0.3 0.54 0.36 0.54 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 12.2442245 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.165 0.895 5.035 0.895 5.035 0.875 5.025 0.875 5.025 0.815 5.085 0.815 5.085 0.56 4.56 0.56 4.56 0.67 4.44 0.67 4.44 0.56 4.255 0.56 4.255 0.88 4.195 0.88 4.195 0.5 5.145 0.5 5.145 0.815 5.165 0.815 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.925 0.975 4.66 0.975 4.66 0.785 4.845 0.785 4.845 0.66 4.925 0.66 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.935 0.805 3.855 0.805 3.855 0.73 3.66 0.73 3.66 0.5 3.74 0.5 3.74 0.645 3.935 0.645 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.815 1.02 0.54 1.02 0.54 1.115 0.46 1.115 0.46 0.94 0.635 0.94 0.635 0.89 0.815 0.89 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 1.77 0 1.77 0 1.65 0.095 1.65 0.095 1.02 0.155 1.02 0.155 1.65 0.505 1.65 0.505 1.215 0.565 1.215 0.565 1.65 1.34 1.65 1.34 1.28 1.4 1.28 1.4 1.65 2.615 1.65 2.615 1.28 2.735 1.28 2.735 1.34 2.675 1.34 2.675 1.65 3.875 1.65 3.875 1.065 3.935 1.065 3.935 1.65 4.675 1.65 4.675 1.25 4.735 1.25 4.735 1.65 5.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 0.06 4.795 0.06 4.795 0.4 4.735 0.4 4.735 0.06 3.935 0.06 3.935 0.4 3.875 0.4 3.875 0.06 2.735 0.06 2.735 0.25 2.615 0.25 2.615 0.19 2.675 0.19 2.675 0.06 1.425 0.06 1.425 0.445 1.365 0.445 1.365 0.06 0.565 0.06 0.565 0.52 0.505 0.52 0.505 0.06 0.155 0.06 0.155 0.52 0.095 0.52 0.095 0.06 0 0.06 0 -0.06 5.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.325 1.135 5.19 1.135 5.19 1.195 5.13 1.195 5.13 1.135 4.43 1.135 4.43 0.82 4.49 0.82 4.49 1.075 5.265 1.075 5.265 0.715 5.245 0.715 5.245 0.42 5.305 0.42 5.305 0.655 5.325 0.655 ;
      POLYGON 4.48 0.4 4.095 0.4 4.095 0.98 4.33 0.98 4.33 1.37 4.27 1.37 4.27 1.04 4.035 1.04 4.035 0.965 3.5 0.965 3.5 1.04 3.44 1.04 3.44 0.44 3.56 0.44 3.56 0.5 3.5 0.5 3.5 0.905 4.035 0.905 4.035 0.34 4.42 0.34 4.42 0.28 4.48 0.28 ;
      POLYGON 3.73 0.4 3.67 0.4 3.67 0.34 3.34 0.34 3.34 1.185 3.73 1.185 3.73 1.245 3.28 1.245 3.28 0.34 2.96 0.34 2.96 0.6 3.02 0.6 3.02 0.66 2.9 0.66 2.9 0.41 2.455 0.41 2.455 0.34 2.135 0.34 2.135 0.645 2.07 0.645 2.07 0.765 1.785 0.765 1.785 0.825 1.725 0.825 1.725 0.705 2.01 0.705 2.01 0.585 2.075 0.585 2.075 0.28 2.515 0.28 2.515 0.35 2.9 0.35 2.9 0.28 3.73 0.28 ;
      POLYGON 3.18 1.18 3.12 1.18 3.12 0.82 2.51 0.82 2.51 0.76 3.12 0.76 3.12 0.5 3.06 0.5 3.06 0.44 3.18 0.44 ;
      POLYGON 3.07 1.34 2.95 1.34 2.95 1.18 2.25 1.18 2.25 1.205 1.63 1.205 1.63 1.18 0.77 1.18 0.77 1.24 0.71 1.24 0.71 1.12 0.915 1.12 0.915 0.54 0.975 0.54 0.975 1.12 1.69 1.12 1.69 1.145 2.19 1.145 2.19 0.74 2.25 0.74 2.25 1.12 3.01 1.12 3.01 1.28 3.07 1.28 ;
      POLYGON 2.8 0.66 2.41 0.66 2.41 1.02 2.35 1.02 2.35 0.57 2.235 0.57 2.235 0.44 2.355 0.44 2.355 0.51 2.41 0.51 2.41 0.6 2.8 0.6 ;
      POLYGON 1.975 0.485 1.91 0.485 1.91 0.605 1.625 0.605 1.625 0.925 1.85 0.925 1.85 1.045 1.79 1.045 1.79 0.985 1.245 0.985 1.245 0.84 1.235 0.84 1.235 0.72 1.305 0.72 1.305 0.925 1.565 0.925 1.565 0.545 1.85 0.545 1.85 0.425 1.975 0.425 ;
      POLYGON 1.465 0.82 1.405 0.82 1.405 0.605 1.135 0.605 1.135 0.9 1.145 0.9 1.145 1.02 1.085 1.02 1.085 0.94 1.075 0.94 1.075 0.44 0.815 0.44 0.815 0.79 0.46 0.79 0.46 0.73 0.755 0.73 0.755 0.38 1.22 0.38 1.22 0.545 1.465 0.545 ;
  END
END SDFFHQX2

MACRO SDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFHQX4 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.60066 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.165 0.715 4.56 0.715 4.56 0.87 4.53 0.87 4.53 0.93 4.47 0.93 4.47 0.81 4.5 0.81 4.5 0.655 5.035 0.655 5.035 0.625 5.165 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.20512825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.82 0.815 5.06 0.985 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.21 0.93 4.13 0.93 4.13 0.92 3.86 0.92 3.86 0.79 3.94 0.79 3.94 0.84 4.13 0.84 4.13 0.75 4.21 0.75 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.69 0.34 1.19 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8383 LAYER Metal1 ;
    ANTENNADIFFAREA 3.66465 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.371025 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.64988875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 60.0283 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.065 1.075 0.46 1.075 0.46 0.79 0.525 0.79 0.525 0.54 0.585 0.54 0.585 0.85 0.54 0.85 0.54 1.015 1.005 1.015 1.005 0.54 1.065 0.54 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 1.77 0 1.77 0 1.65 0.27 1.65 0.27 1.51 0.33 1.51 0.33 1.65 0.71 1.65 0.71 1.45 0.83 1.45 0.83 1.51 0.77 1.51 0.77 1.65 1.18 1.65 1.18 1.45 1.3 1.45 1.3 1.51 1.24 1.51 1.24 1.65 1.65 1.65 1.65 1.45 1.77 1.45 1.77 1.51 1.71 1.51 1.71 1.65 2.85 1.65 2.85 1.4 2.97 1.4 2.97 1.46 2.91 1.46 2.91 1.65 4.19 1.65 4.19 1.26 4.25 1.26 4.25 1.65 4.915 1.65 4.915 1.26 4.975 1.26 4.975 1.65 5.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 0.06 5.05 0.06 5.05 0.525 4.99 0.525 4.99 0.06 4.18 0.06 4.18 0.55 4.12 0.55 4.12 0.06 2.97 0.06 2.97 0.255 2.85 0.255 2.85 0.195 2.91 0.195 2.91 0.06 1.71 0.06 1.71 0.52 1.65 0.52 1.65 0.06 1.29 0.06 1.29 0.52 1.23 0.52 1.23 0.06 0.79 0.06 0.79 0.52 0.73 0.52 0.73 0.06 0.38 0.06 0.38 0.52 0.32 0.52 0.32 0.06 0 0.06 0 -0.06 5.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.325 1.145 5.255 1.145 5.255 1.205 5.195 1.205 5.195 1.145 4.66 1.145 4.66 0.83 4.72 0.83 4.72 1.085 5.265 1.085 5.265 0.43 5.325 0.43 ;
      POLYGON 4.74 0.555 4.4 0.555 4.4 0.71 4.37 0.71 4.37 1.03 4.56 1.03 4.56 1.38 4.5 1.38 4.5 1.09 3.625 1.09 3.625 1.03 3.685 1.03 3.685 0.515 3.805 0.515 3.805 0.575 3.745 0.575 3.745 1.03 4.31 1.03 4.31 0.65 4.34 0.65 4.34 0.495 4.68 0.495 4.68 0.435 4.74 0.435 ;
      POLYGON 4.075 1.255 3.465 1.255 3.465 0.81 3.525 0.81 3.525 0.415 3.205 0.415 3.205 0.775 3.145 0.775 3.145 0.415 2.37 0.415 2.37 0.725 2.335 0.725 2.335 0.785 2.07 0.785 2.07 0.905 2.01 0.905 2.01 0.725 2.275 0.725 2.275 0.665 2.31 0.665 2.31 0.355 3.975 0.355 3.975 0.55 3.915 0.55 3.915 0.415 3.585 0.415 3.585 0.93 3.525 0.93 3.525 1.195 4.075 1.195 ;
      POLYGON 3.425 0.575 3.365 0.575 3.365 1.265 3.305 1.265 3.305 0.935 2.765 0.935 2.765 0.845 2.885 0.845 2.885 0.875 3.305 0.875 3.305 0.515 3.425 0.515 ;
      POLYGON 3.255 1.425 3.135 1.425 3.135 1.3 2.505 1.3 2.505 1.35 0.085 1.35 0.085 0.54 0.145 0.54 0.145 1.29 2.445 1.29 2.445 0.8 2.505 0.8 2.505 1.24 3.195 1.24 3.195 1.365 3.255 1.365 ;
      POLYGON 3.045 0.745 2.665 0.745 2.665 1.14 2.605 1.14 2.605 0.575 2.47 0.575 2.47 0.515 2.665 0.515 2.665 0.685 3.045 0.685 ;
      POLYGON 2.21 0.565 1.91 0.565 1.91 1.005 2.145 1.005 2.145 1.19 2.085 1.19 2.085 1.065 1.85 1.065 1.85 0.925 1.52 0.925 1.52 0.805 1.58 0.805 1.58 0.865 1.85 0.865 1.85 0.505 2.21 0.505 ;
      POLYGON 1.75 0.765 1.69 0.765 1.69 0.705 1.42 0.705 1.42 1.025 1.535 1.025 1.535 1.085 1.36 1.085 1.36 0.705 1.225 0.705 1.225 0.82 1.165 0.82 1.165 0.645 1.445 0.645 1.445 0.485 1.505 0.485 1.505 0.645 1.75 0.645 ;
  END
END SDFFHQX4

MACRO SDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFHQX8 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.21782175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 0.745 6.34 0.745 6.34 0.705 5.685 0.705 5.685 0.755 5.595 0.755 5.595 0.965 5.535 0.965 5.535 0.695 5.625 0.695 5.625 0.645 6.235 0.645 6.235 0.625 6.4 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.24 0.885 6.165 0.885 6.165 1.01 5.865 1.01 5.865 0.805 6.24 0.805 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.275 1.015 5.195 1.015 5.195 0.92 5.06 0.92 5.06 0.65 5.14 0.65 5.14 0.79 5.275 0.79 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.83 0.895 2.555 0.895 2.555 0.815 2.72 0.815 2.72 0.59 2.83 0.59 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6952 LAYER Metal1 ;
    ANTENNADIFFAREA 4.57105 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.528525 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.991533 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 54.8034625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.36 0.65 1.315 0.65 1.315 0.9 1.36 0.9 1.36 1.345 1.3 1.345 1.3 0.96 1.255 0.96 1.255 0.8 0.95 0.8 0.95 1.345 0.89 1.345 0.89 0.73 0.54 0.73 0.54 1.345 0.48 1.345 0.48 0.73 0.13 0.73 0.13 1.345 0.07 1.345 0.07 0.73 0.06 0.73 0.06 0.6 0.07 0.6 0.07 0.54 0.14 0.54 0.14 0.67 0.48 0.67 0.48 0.54 0.54 0.54 0.54 0.67 0.89 0.67 0.89 0.54 0.95 0.54 0.95 0.74 1.255 0.74 1.255 0.59 1.3 0.59 1.3 0.53 1.36 0.53 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 1.77 0 1.77 0 1.65 0.275 1.65 0.275 0.9 0.335 0.9 0.335 1.65 0.685 1.65 0.685 0.9 0.745 0.9 0.745 1.65 1.095 1.65 1.095 0.9 1.155 0.9 1.155 1.65 1.505 1.65 1.505 0.905 1.565 0.905 1.565 1.65 1.945 1.65 1.945 1.055 2.005 1.055 2.005 1.65 2.93 1.65 2.93 1.51 2.99 1.51 2.99 1.65 4.055 1.65 4.055 1.315 4.175 1.315 4.175 1.375 4.115 1.375 4.115 1.65 5.235 1.65 5.235 1.285 5.295 1.285 5.295 1.65 6.055 1.65 6.055 1.285 6.115 1.285 6.115 1.65 6.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 0.06 6.115 0.06 6.115 0.525 6.055 0.525 6.055 0.06 5.365 0.06 5.365 0.435 5.305 0.435 5.305 0.06 4.175 0.06 4.175 0.17 4.055 0.17 4.055 0.06 2.915 0.06 2.915 0.17 2.795 0.17 2.795 0.06 1.975 0.06 1.975 0.485 1.915 0.485 1.915 0.06 1.565 0.06 1.565 0.485 1.505 0.485 1.505 0.06 1.155 0.06 1.155 0.485 1.095 0.485 1.095 0.06 0.745 0.06 0.745 0.485 0.685 0.485 0.685 0.06 0.335 0.06 0.335 0.485 0.275 0.485 0.275 0.06 0 0.06 0 -0.06 6.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.56 1.17 6.35 1.17 6.35 1.23 6.29 1.23 6.29 1.17 5.705 1.17 5.705 0.855 5.765 0.855 5.765 1.11 6.5 1.11 6.5 0.525 6.29 0.525 6.29 0.405 6.35 0.405 6.35 0.465 6.56 0.465 ;
      POLYGON 5.805 0.545 5.525 0.545 5.525 0.595 5.435 0.595 5.435 1.115 5.605 1.115 5.605 1.405 5.545 1.405 5.545 1.175 4.84 1.175 4.84 0.98 4.9 0.98 4.9 0.515 4.84 0.515 4.84 0.455 4.96 0.455 4.96 1.115 5.375 1.115 5.375 0.535 5.465 0.535 5.465 0.485 5.745 0.485 5.745 0.425 5.805 0.425 ;
      POLYGON 5.13 0.55 5.07 0.55 5.07 0.355 4.74 0.355 4.74 1.315 5.12 1.315 5.12 1.375 4.68 1.375 4.68 0.355 4.36 0.355 4.36 0.615 4.41 0.615 4.41 0.735 4.3 0.735 4.3 0.355 3.575 0.355 3.575 0.615 3.69 0.615 3.69 0.735 3.63 0.735 3.63 0.675 3.515 0.675 3.515 0.295 5.13 0.295 ;
      POLYGON 4.58 1.215 4.52 1.215 4.52 0.895 4.01 0.895 4.01 0.855 3.95 0.855 3.95 0.795 4.07 0.795 4.07 0.835 4.52 0.835 4.52 0.515 4.46 0.515 4.46 0.455 4.58 0.455 ;
      POLYGON 4.47 1.375 4.35 1.375 4.35 1.215 3.09 1.215 3.09 0.49 2.455 0.49 2.455 0.995 2.705 0.995 2.705 1.115 2.645 1.115 2.645 1.055 2.395 1.055 2.395 0.43 3.15 0.43 3.15 1.155 3.47 1.155 3.47 0.835 3.41 0.835 3.41 0.775 3.53 0.775 3.53 1.155 4.41 1.155 4.41 1.315 4.47 1.315 ;
      POLYGON 4.2 0.715 4.14 0.715 4.14 0.695 3.85 0.695 3.85 1.055 3.79 1.055 3.79 0.515 3.675 0.515 3.675 0.455 3.85 0.455 3.85 0.635 4.14 0.635 4.14 0.595 4.2 0.595 ;
      POLYGON 3.37 1.055 3.31 1.055 3.31 0.995 3.25 0.995 3.25 0.33 2.135 0.33 2.135 0.795 2.075 0.795 2.075 0.27 3.31 0.27 3.31 0.935 3.37 0.935 ;
      POLYGON 2.99 1.275 2.21 1.275 2.21 1.345 2.15 1.345 2.15 0.955 1.8 0.955 1.8 1.345 1.74 1.345 1.74 0.955 1.71 0.955 1.71 0.805 1.415 0.805 1.415 0.745 1.71 0.745 1.71 0.505 1.77 0.505 1.77 0.895 2.235 0.895 2.235 0.505 2.295 0.505 2.295 1.215 2.93 1.215 2.93 0.74 2.99 0.74 ;
  END
END SDFFHQX8

MACRO SDFFNSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSRX1 0 0 ;
  SIZE 7.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3272 LAYER Metal1 ;
    ANTENNADIFFAREA 4.1535 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2691 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.0802675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 124.45930875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 0.635 0.95 0.635 0.95 1.035 0.995 1.035 0.995 1.425 0.935 1.425 0.935 1.11 0.86 1.11 0.86 0.98 0.89 0.98 0.89 0.555 0.94 0.555 0.94 0.515 1 0.515 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3272 LAYER Metal1 ;
    ANTENNADIFFAREA 4.1535 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2691 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.0802675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 124.45930875 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.325 1.29 0.245 1.29 0.245 0.73 0.06 0.73 0.06 0.6 0.245 0.6 0.245 0.54 0.325 0.54 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.52 0.725 7.04 0.725 7.04 0.645 7.235 0.645 7.235 0.625 7.365 0.625 7.365 0.645 7.52 0.645 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.2 0.825 7.52 1.085 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.56 1.15 6.46 1.15 6.46 0.98 6.48 0.98 6.48 0.67 6.56 0.67 ;
    END
  END D
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.36 1.15 6.28 1.15 6.28 0.92 6.26 0.92 6.26 0.67 6.36 0.67 ;
    END
  END CKN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 27.54629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.515 1.405 4.06 1.405 4.06 1.235 3.16 1.235 3.16 0.985 2.305 0.985 2.305 0.895 2.13 0.895 2.13 0.835 2.235 0.835 2.235 0.815 2.365 0.815 2.365 0.925 3.22 0.925 3.22 1.175 4.12 1.175 4.12 1.345 4.515 1.345 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 1.205 1.095 1.205 1.095 1.005 1.245 1.005 1.245 0.895 1.365 0.895 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.8 1.77 0 1.77 0 1.65 0.47 1.65 0.47 0.995 0.53 0.995 0.53 1.65 1.14 1.65 1.14 1.305 1.2 1.305 1.2 1.65 1.985 1.65 1.985 1.155 2.045 1.155 2.045 1.65 2.74 1.65 2.74 1.425 2.86 1.425 2.86 1.485 2.8 1.485 2.8 1.65 3.67 1.65 3.67 1.54 3.79 1.54 3.79 1.65 4.615 1.65 4.615 1.49 4.735 1.49 4.735 1.55 4.675 1.55 4.675 1.65 5.825 1.65 5.825 0.995 5.885 0.995 5.885 1.65 6.44 1.65 6.44 1.25 6.5 1.25 6.5 1.65 7.285 1.65 7.285 1.345 7.405 1.345 7.405 1.405 7.345 1.405 7.345 1.65 7.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.8 0.06 7.36 0.06 7.36 0.44 7.3 0.44 7.3 0.06 6.535 0.06 6.535 0.41 6.415 0.41 6.415 0.35 6.475 0.35 6.475 0.06 5.775 0.06 5.775 0.17 5.655 0.17 5.655 0.06 4.675 0.06 4.675 0.56 4.615 0.56 4.615 0.06 2.015 0.06 2.015 0.2 1.955 0.2 1.955 0.06 1.205 0.06 1.205 0.635 1.145 0.635 1.145 0.06 0.53 0.06 0.53 0.635 0.47 0.635 0.47 0.06 0 0.06 0 -0.06 7.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.68 1.245 7.58 1.245 7.58 1.34 7.52 1.34 7.52 1.245 7.1 1.245 7.1 1.405 6.66 1.405 6.66 0.675 6.78 0.675 6.78 0.735 6.72 0.735 6.72 1.345 7.04 1.345 7.04 0.995 7.1 0.995 7.1 1.185 7.62 1.185 7.62 0.465 7.505 0.465 7.505 0.345 7.565 0.345 7.565 0.405 7.68 0.405 ;
      POLYGON 6.94 1.245 6.82 1.245 6.82 0.835 6.88 0.835 6.88 0.57 6.255 0.57 6.255 0.37 5.935 0.37 5.935 0.4 5.3 0.4 5.3 0.5 5.52 0.5 5.52 0.88 5.46 0.88 5.46 1.11 5.4 1.11 5.4 0.82 5.46 0.82 5.46 0.56 5.24 0.56 5.24 0.34 5.875 0.34 5.875 0.31 6.315 0.31 6.315 0.51 6.755 0.51 6.755 0.345 6.815 0.345 6.815 0.51 6.94 0.51 ;
      POLYGON 6.295 1.37 6.235 1.37 6.235 1.31 6.035 1.31 6.035 0.785 5.84 0.785 5.84 0.845 5.78 0.845 5.78 0.725 6.035 0.725 6.035 0.47 6.155 0.47 6.155 0.53 6.095 0.53 6.095 1.25 6.295 1.25 ;
      POLYGON 5.74 0.625 5.68 0.625 5.68 1.335 4.86 1.335 4.86 1.245 4.22 1.245 4.22 1.075 3.885 1.075 3.885 0.83 3.945 0.83 3.945 1.015 4.28 1.015 4.28 1.185 4.86 1.185 4.86 0.895 4.98 0.895 4.98 1.015 4.92 1.015 4.92 1.275 5.24 1.275 5.24 0.66 5.36 0.66 5.36 0.72 5.3 0.72 5.3 1.275 5.62 1.275 5.62 0.565 5.74 0.565 ;
      POLYGON 5.14 1.175 5.02 1.175 5.02 1.115 5.08 1.115 5.08 0.755 4.32 0.755 4.32 0.635 4.38 0.635 4.38 0.695 5.08 0.695 5.08 0.585 5.035 0.585 5.035 0.465 5.095 0.465 5.095 0.525 5.14 0.525 ;
      POLYGON 4.76 0.915 4.44 0.915 4.44 1.025 4.5 1.025 4.5 1.085 4.38 1.085 4.38 0.915 4.16 0.915 4.16 0.69 3.785 0.69 3.785 1.055 3.54 1.055 3.54 0.995 3.725 0.995 3.725 0.66 3.64 0.66 3.64 0.54 3.7 0.54 3.7 0.6 3.785 0.6 3.785 0.63 4.16 0.63 4.16 0.465 4.22 0.465 4.22 0.855 4.76 0.855 ;
      POLYGON 4.485 0.53 4.32 0.53 4.32 0.365 4.045 0.365 4.045 0.53 3.925 0.53 3.925 0.47 3.985 0.47 3.985 0.305 4.38 0.305 4.38 0.47 4.485 0.47 ;
      POLYGON 3.96 1.395 2.96 1.395 2.96 1.325 2.64 1.325 2.64 1.485 2.52 1.485 2.52 1.365 2.145 1.365 2.145 1.055 1.885 1.055 1.885 1.34 1.465 1.34 1.465 0.54 1.525 0.54 1.525 1.28 1.825 1.28 1.825 0.995 2.205 0.995 2.205 1.305 2.58 1.305 2.58 1.265 3.02 1.265 3.02 1.335 3.96 1.335 ;
      POLYGON 3.625 0.895 3.565 0.895 3.565 0.835 3.48 0.835 3.48 0.265 3.225 0.265 3.225 0.205 3.54 0.205 3.54 0.775 3.625 0.775 ;
      POLYGON 3.44 1.05 3.32 1.05 3.32 0.825 2.465 0.825 2.465 0.715 1.97 0.715 1.97 0.775 1.91 0.775 1.91 0.655 2.525 0.655 2.525 0.765 3.32 0.765 3.32 0.54 3.38 0.54 3.38 0.99 3.44 0.99 ;
      POLYGON 3.175 0.665 2.625 0.665 2.625 0.42 2.705 0.42 2.705 0.585 3.095 0.585 3.095 0.54 3.175 0.54 ;
      POLYGON 3.06 1.165 2.385 1.165 2.385 1.205 2.305 1.205 2.305 1.085 3.06 1.085 ;
      POLYGON 2.925 0.485 2.805 0.485 2.805 0.32 2.525 0.32 2.525 0.485 2.275 0.485 2.275 0.425 2.465 0.425 2.465 0.26 2.865 0.26 2.865 0.425 2.925 0.425 ;
      POLYGON 2.365 0.325 2.175 0.325 2.175 0.555 1.835 0.555 1.835 0.58 1.725 0.58 1.725 1.18 1.665 1.18 1.665 0.52 1.78 0.52 1.78 0.42 1.365 0.42 1.365 0.795 1.05 0.795 1.05 0.735 1.305 0.735 1.305 0.36 1.84 0.36 1.84 0.495 2.115 0.495 2.115 0.265 2.365 0.265 ;
      POLYGON 0.76 1.02 0.68 1.02 0.68 0.815 0.425 0.815 0.425 0.735 0.68 0.735 0.68 0.54 0.76 0.54 ;
  END
END SDFFNSRX1

MACRO SDFFNSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSRX2 0 0 ;
  SIZE 8.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.531125 LAYER Metal1 ;
    ANTENNADIFFAREA 4.5961 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.334575 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.5429275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 105.7206905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.02 0.99 7.885 0.99 7.885 0.705 7.835 0.705 7.835 0.625 7.885 0.625 7.885 0.535 7.91 0.535 7.91 0.495 7.99 0.495 7.99 0.615 7.965 0.615 7.965 0.91 8.02 0.91 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.581125 LAYER Metal1 ;
    ANTENNADIFFAREA 4.5961 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.334575 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.692371 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 106.35283575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.465 1.41 7.405 1.41 7.405 1.11 7.26 1.11 7.26 0.98 7.405 0.98 7.405 0.495 7.465 0.495 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.64 0.545 0.56 0.545 0.56 0.54 0.195 0.54 0.195 0.46 0.46 0.46 0.46 0.41 0.54 0.41 0.54 0.42 0.64 0.42 ;
    END
  END SE
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.186 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.74074075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 63.888889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.465 0.705 3.26 0.705 3.26 0.33 3.34 0.33 3.34 0.625 3.465 0.625 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.06 0.65 1.14 1.15 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.46 1.02 0.26 1.02 0.26 0.79 0.38 0.79 0.38 0.64 0.46 0.64 ;
    END
  END SI
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.06 0.69 7.14 1.19 ;
    END
  END RN
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.605 0.895 1.335 0.895 1.335 0.585 1.415 0.585 1.415 0.815 1.605 0.815 ;
    END
  END CKN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.6 1.77 0 1.77 0 1.65 0.285 1.65 0.285 1.51 0.345 1.51 0.345 1.65 1.135 1.65 1.135 1.25 1.195 1.25 1.195 1.65 2.21 1.65 2.21 1.04 2.33 1.04 2.33 1.1 2.27 1.1 2.27 1.65 3.375 1.65 3.375 1.285 3.435 1.285 3.435 1.65 4.235 1.65 4.235 1.415 4.355 1.415 4.355 1.475 4.295 1.475 4.295 1.65 5.71 1.65 5.71 1.385 5.77 1.385 5.77 1.65 6.55 1.65 6.55 1.51 6.61 1.51 6.61 1.65 7.2 1.65 7.2 1.29 7.26 1.29 7.26 1.65 7.61 1.65 7.61 1.32 7.73 1.32 7.73 1.38 7.67 1.38 7.67 1.65 8.15 1.65 8.15 1.25 8.27 1.25 8.27 1.31 8.21 1.31 8.21 1.65 8.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.6 0.06 8.195 0.06 8.195 0.59 8.135 0.59 8.135 0.06 7.785 0.06 7.785 0.475 7.725 0.475 7.725 0.06 7.26 0.06 7.26 0.17 7.14 0.17 7.14 0.06 6.57 0.06 6.57 0.575 6.51 0.575 6.51 0.06 3.785 0.06 3.785 0.535 3.725 0.535 3.725 0.06 2.195 0.06 2.195 0.17 2.075 0.17 2.075 0.06 1.34 0.06 1.34 0.325 1.22 0.325 1.22 0.265 1.28 0.265 1.28 0.06 0.36 0.06 0.36 0.355 0.3 0.355 0.3 0.06 0 0.06 0 -0.06 8.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 8.475 1.245 8.415 1.245 8.415 0.775 8.065 0.775 8.065 0.715 8.34 0.715 8.34 0.495 8.4 0.495 8.4 0.715 8.475 0.715 ;
      POLYGON 8.315 1.15 7.565 1.15 7.565 0.37 7.305 0.37 7.305 0.785 7.245 0.785 7.245 0.37 6.775 0.37 6.775 0.675 6.8 0.675 6.8 1.015 6.78 1.015 6.78 1.085 6.72 1.085 6.72 0.965 6.74 0.965 6.74 0.735 6.3 0.735 6.3 0.795 6.24 0.795 6.24 0.675 6.715 0.675 6.715 0.31 7.625 0.31 7.625 1.09 8.255 1.09 8.255 0.955 8.315 0.955 ;
      POLYGON 7.055 0.59 6.96 0.59 6.96 1.29 7.055 1.29 7.055 1.41 6.56 1.41 6.56 1.275 6.03 1.275 6.03 1.215 6.62 1.215 6.62 1.35 6.9 1.35 6.9 0.53 6.995 0.53 6.995 0.47 7.055 0.47 ;
      POLYGON 6.64 0.895 6.46 0.895 6.46 0.955 5.215 0.955 5.215 1.05 5.155 1.05 5.155 0.51 5.275 0.51 5.275 0.57 5.215 0.57 5.215 0.895 6.4 0.895 6.4 0.835 6.64 0.835 ;
      POLYGON 6.46 1.435 5.87 1.435 5.87 1.285 5.61 1.285 5.61 1.34 4.455 1.34 4.455 1.315 4.135 1.315 4.135 1.345 3.62 1.345 3.62 1.285 4.075 1.285 4.075 1.255 4.515 1.255 4.515 1.28 5.55 1.28 5.55 1.225 5.93 1.225 5.93 1.375 6.46 1.375 ;
      RECT 5.33 1.055 6.395 1.115 ;
      POLYGON 6.37 0.575 6.29 0.575 6.29 0.41 5.97 0.41 5.97 0.575 5.89 0.575 5.89 0.33 6.37 0.33 ;
      POLYGON 6.19 0.57 6.13 0.57 6.13 0.735 5.39 0.735 5.39 0.48 5.45 0.48 5.45 0.675 6.07 0.675 6.07 0.51 6.19 0.51 ;
      POLYGON 5.34 0.235 5.055 0.235 5.055 1.18 4.615 1.18 4.615 1.155 3.975 1.155 3.975 1.185 3.18 1.185 3.18 1.315 3.06 1.315 3.06 1.185 2.445 1.185 2.445 0.9 2.455 0.9 2.455 0.545 2.575 0.545 2.575 0.605 2.515 0.605 2.515 0.96 2.505 0.96 2.505 1.125 2.835 1.125 2.835 0.635 2.895 0.635 2.895 1.125 3.915 1.125 3.915 1.095 4.675 1.095 4.675 1.12 4.995 1.12 4.995 0.175 5.34 0.175 ;
      POLYGON 4.895 1.02 4.775 1.02 4.775 0.96 4.835 0.96 4.835 0.86 3.755 0.86 3.755 0.965 3.815 0.965 3.815 1.025 3.695 1.025 3.695 0.865 3.24 0.865 3.24 0.805 3.72 0.805 3.72 0.8 4.15 0.8 4.15 0.44 4.21 0.44 4.21 0.8 4.835 0.8 4.835 0.48 4.895 0.48 ;
      POLYGON 4.415 0.535 4.355 0.535 4.355 0.34 3.99 0.34 3.99 0.535 3.93 0.535 3.93 0.28 4.415 0.28 ;
      POLYGON 4.05 0.7 3.565 0.7 3.565 0.23 3.115 0.23 3.115 1.025 2.995 1.025 2.995 0.965 3.055 0.965 3.055 0.505 2.995 0.505 2.995 0.445 3.055 0.445 3.055 0.17 3.625 0.17 3.625 0.64 4.05 0.64 ;
      POLYGON 2.82 0.535 2.735 0.535 2.735 1.025 2.615 1.025 2.615 0.965 2.675 0.965 2.675 0.475 2.76 0.475 2.76 0.375 2.355 0.375 2.355 0.47 1.5 0.47 1.5 0.485 0.8 0.485 0.8 1.34 0.605 1.34 0.605 1.28 0.74 1.28 0.74 0.26 0.8 0.26 0.8 0.425 1.44 0.425 1.44 0.41 2.295 0.41 2.295 0.315 2.82 0.315 ;
      POLYGON 2.355 0.8 1.765 0.8 1.765 1.245 1.4 1.245 1.4 1.185 1.705 1.185 1.705 0.63 1.6 0.63 1.6 0.57 1.765 0.57 1.765 0.74 2.355 0.74 ;
      POLYGON 0.96 1.5 0.445 1.5 0.445 1.18 0.155 1.18 0.155 1.24 0.095 1.24 0.095 1.18 0.035 1.18 0.035 0.295 0.09 0.295 0.09 0.235 0.15 0.235 0.15 0.355 0.095 0.355 0.095 1.12 0.56 1.12 0.56 0.995 0.62 0.995 0.62 1.18 0.505 1.18 0.505 1.44 0.9 1.44 0.9 0.6 0.96 0.6 ;
  END
END SDFFNSRX2

MACRO SDFFNSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSRX4 0 0 ;
  SIZE 9.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.308375 LAYER Metal1 ;
    ANTENNADIFFAREA 5.4387 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4878 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.8822775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 85.0553505 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.67 0.54 8.14 0.54 8.14 0.915 8.515 0.915 8.515 1.305 8.455 1.305 8.455 0.975 8.105 0.975 8.105 1.305 8.045 1.305 8.045 0.915 8.06 0.915 8.06 0.79 8.08 0.79 8.08 0.48 8.67 0.48 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.308375 LAYER Metal1 ;
    ANTENNADIFFAREA 5.4387 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4878 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.8822775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 85.0553505 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.73 0.54 7.32 0.54 7.32 0.79 7.34 0.79 7.34 0.86 7.695 0.86 7.695 1.305 7.635 1.305 7.635 0.92 7.32 0.92 7.32 1.305 7.225 1.305 7.225 0.915 7.26 0.915 7.26 0.54 7.14 0.54 7.14 0.48 7.73 0.48 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 12.31481475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.59 0.735 4.085 0.735 4.085 0.705 4.035 0.705 4.035 0.625 4.165 0.625 4.165 0.655 4.59 0.655 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.935 0.905 3.855 0.905 3.855 0.705 3.635 0.705 3.635 0.625 3.935 0.625 ;
    END
  END SN
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.7 1.54 1.2 ;
    END
  END CKN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.65 1.34 1.15 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.68 0.92 0.54 0.92 0.54 1.075 0.46 1.075 0.46 0.715 0.68 0.715 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 19.675926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.16 1.06 1.1 1.06 1.1 0.355 0.84 0.355 0.84 0.795 0.78 0.795 0.78 0.615 0.36 0.615 0.36 0.675 0.3 0.675 0.3 0.555 0.66 0.555 0.66 0.41 0.78 0.41 0.78 0.295 1.16 0.295 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.4 1.77 0 1.77 0 1.65 0.535 1.65 0.535 1.335 0.595 1.335 0.595 1.65 1.365 1.65 1.365 1.51 1.425 1.51 1.425 1.65 2.595 1.65 2.595 1.55 2.535 1.55 2.535 1.49 2.655 1.49 2.655 1.65 2.995 1.65 2.995 1.54 3.115 1.54 3.115 1.65 3.93 1.65 3.93 1.49 4.05 1.49 4.05 1.55 3.99 1.55 3.99 1.65 5.865 1.65 5.865 1.215 5.985 1.215 5.985 1.275 5.925 1.275 5.925 1.65 6.41 1.65 6.41 1.185 6.47 1.185 6.47 1.65 6.935 1.65 6.935 0.995 6.995 0.995 6.995 1.65 7.43 1.65 7.43 1.02 7.49 1.02 7.49 1.65 7.84 1.65 7.84 0.915 7.9 0.915 7.9 1.65 8.25 1.65 8.25 1.075 8.31 1.075 8.31 1.65 8.685 1.65 8.685 0.96 8.745 0.96 8.745 1.65 9.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.4 0.06 8.99 0.06 8.99 0.43 8.93 0.43 8.93 0.06 8.435 0.06 8.435 0.17 8.315 0.17 8.315 0.06 7.965 0.06 7.965 0.17 7.845 0.17 7.845 0.06 7.495 0.06 7.495 0.17 7.375 0.17 7.375 0.06 6.88 0.06 6.88 0.485 6.82 0.485 6.82 0.06 6.47 0.06 6.47 0.485 6.41 0.485 6.41 0.06 4.545 0.06 4.545 0.395 4.425 0.395 4.425 0.335 4.485 0.335 4.485 0.06 2.78 0.06 2.78 0.17 2.66 0.17 2.66 0.06 1.36 0.06 1.36 0.55 1.3 0.55 1.3 0.06 0.435 0.06 0.435 0.455 0.375 0.455 0.375 0.06 0 0.06 0 -0.06 9.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 9.195 0.86 8.95 0.86 8.95 1.305 8.89 1.305 8.89 0.86 8.615 0.86 8.615 0.71 8.735 0.71 8.735 0.8 9.135 0.8 9.135 0.45 9.195 0.45 ;
      POLYGON 9.035 0.7 8.835 0.7 8.835 0.59 8.77 0.59 8.77 0.38 7.04 0.38 7.04 0.645 6.79 0.645 6.79 0.745 7.12 0.745 7.12 0.805 6.79 0.805 6.79 1.305 6.73 1.305 6.73 0.66 6.1 0.66 6.1 0.6 6.615 0.6 6.615 0.45 6.675 0.45 6.675 0.585 6.98 0.585 6.98 0.32 8.83 0.32 8.83 0.53 8.895 0.53 8.895 0.64 9.035 0.64 ;
      POLYGON 6.63 0.955 5.24 0.955 5.24 1.145 5.18 1.145 5.18 0.66 5.16 0.66 5.16 0.54 5.22 0.54 5.22 0.61 5.24 0.61 5.24 0.895 6.51 0.895 6.51 0.855 6.63 0.855 ;
      POLYGON 6.295 1.18 6.085 1.18 6.085 1.115 5.355 1.115 5.355 1.055 6.145 1.055 6.145 1.12 6.295 1.12 ;
      POLYGON 6.265 0.485 6.185 0.485 6.185 0.32 5.82 0.32 5.82 0.455 5.7 0.455 5.7 0.375 5.74 0.375 5.74 0.24 6.265 0.24 ;
      POLYGON 6.085 0.5 6 0.5 6 0.635 5.5 0.635 5.5 0.515 5.58 0.515 5.58 0.555 5.92 0.555 5.92 0.42 6.085 0.42 ;
      POLYGON 5.955 0.795 5.34 0.795 5.34 0.415 4.75 0.415 4.75 0.99 4.63 0.99 4.63 0.93 4.69 0.93 4.69 0.555 4.265 0.555 4.265 0.29 3.96 0.29 3.96 0.23 4.325 0.23 4.325 0.495 4.69 0.495 4.69 0.355 5.4 0.355 5.4 0.735 5.955 0.735 ;
      POLYGON 5.645 1.34 5.525 1.34 5.525 1.31 4.31 1.31 4.31 1.225 3.535 1.225 3.535 1.025 2.995 1.025 2.995 0.9 3.055 0.9 3.055 0.965 3.595 0.965 3.595 1.165 4.37 1.165 4.37 1.25 5.02 1.25 5.02 0.735 5.08 0.735 5.08 1.25 5.585 1.25 5.585 1.28 5.645 1.28 ;
      POLYGON 5.14 1.47 4.15 1.47 4.15 1.385 3.375 1.385 3.375 1.185 2.77 1.185 2.77 1.125 2.835 1.125 2.835 0.99 2.34 0.99 2.34 1.05 2.28 1.05 2.28 0.93 2.835 0.93 2.835 0.63 2.775 0.63 2.775 0.57 2.895 0.57 2.895 1.125 3.435 1.125 3.435 1.325 4.21 1.325 4.21 1.41 5.14 1.41 ;
      POLYGON 5.015 0.635 4.92 0.635 4.92 1.15 4.47 1.15 4.47 1.065 3.695 1.065 3.695 0.865 3.475 0.865 3.475 0.715 3.135 0.715 3.135 0.47 2.5 0.47 2.5 0.445 2.44 0.445 2.44 0.385 2.56 0.385 2.56 0.41 3.195 0.41 3.195 0.655 3.475 0.655 3.475 0.465 3.68 0.465 3.68 0.525 3.535 0.525 3.535 0.805 3.755 0.805 3.755 1.005 4.53 1.005 4.53 1.09 4.86 1.09 4.86 0.575 4.955 0.575 4.955 0.515 5.015 0.515 ;
      POLYGON 3.9 0.525 3.78 0.525 3.78 0.365 3.375 0.365 3.375 0.555 3.295 0.555 3.295 0.285 3.86 0.285 3.86 0.445 3.9 0.445 ;
      POLYGON 3.745 1.545 3.215 1.545 3.215 1.39 2.12 1.39 2.12 0.54 2.18 0.54 2.18 1.33 3.275 1.33 3.275 1.485 3.745 1.485 ;
      POLYGON 2.735 0.83 2.28 0.83 2.28 0.44 2.02 0.44 2.02 0.96 1.96 0.96 1.96 0.44 1.605 0.44 1.605 0.54 1.7 0.54 1.7 1.195 1.64 1.195 1.64 0.6 1.545 0.6 1.545 0.38 2.34 0.38 2.34 0.71 2.36 0.71 2.36 0.77 2.735 0.77 ;
      POLYGON 1.945 1.36 0.94 1.36 0.94 0.455 1 0.455 1 1.3 1.885 1.3 1.885 1.16 1.8 1.16 1.8 0.54 1.86 0.54 1.86 1.1 1.945 1.1 ;
      POLYGON 0.84 1.235 0.39 1.235 0.39 1.36 0.33 1.36 0.33 1.235 0.14 1.235 0.14 0.36 0.2 0.36 0.2 1.175 0.78 1.175 0.78 1.08 0.84 1.08 ;
  END
END SDFFNSRX4

MACRO SDFFNSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFNSRXL 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.288575 LAYER Metal1 ;
    ANTENNADIFFAREA 4.1863 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.243 LAYER Metal1 ;
      ANTENNAMAXAREACAR 17.64845675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 133.45679 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.175 0.49 1.115 0.49 1.115 1.18 1.175 1.18 1.175 1.3 0.86 1.3 0.86 1.17 1.035 1.17 1.035 0.41 1.095 0.41 1.095 0.37 1.175 0.37 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.288575 LAYER Metal1 ;
    ANTENNADIFFAREA 4.1863 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.243 LAYER Metal1 ;
      ANTENNAMAXAREACAR 17.64845675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 133.45679 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.325 1.02 0.245 1.02 0.245 0.73 0.06 0.73 0.06 0.6 0.245 0.6 0.245 0.54 0.325 0.54 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.41666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.765 0.705 7.705 0.705 7.705 0.745 7.645 0.745 7.645 0.725 7.31 0.725 7.31 0.785 7.145 0.785 7.145 1.05 7.085 1.05 7.085 0.665 7.635 0.665 7.635 0.625 7.765 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.765 1.085 7.635 1.085 7.635 0.935 7.415 0.935 7.415 0.855 7.765 0.855 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.825 1.085 6.515 1.085 6.515 1.005 6.635 1.005 6.635 0.815 6.765 0.815 6.765 1.005 6.825 1.005 ;
    END
  END D
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.415 0.905 6.295 0.905 6.295 1.005 6.415 1.005 6.415 1.085 6.215 1.085 6.215 0.825 6.415 0.825 ;
    END
  END CKN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 28.56481475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.805 1.365 4.35 1.365 4.35 1.235 2.28 1.235 2.28 1.11 2.26 1.11 2.26 0.825 2.32 0.825 2.32 0.98 2.34 0.98 2.34 1.175 4.41 1.175 4.41 1.305 4.805 1.305 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.25925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 0.75 1.565 1.12 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 1.77 0 1.77 0 1.65 0.495 1.65 0.495 0.995 0.555 0.995 0.555 1.65 1.32 1.65 1.32 1.22 1.38 1.22 1.38 1.65 2.22 1.65 2.22 1.54 2.34 1.54 2.34 1.65 2.94 1.65 2.94 1.54 3.06 1.54 3.06 1.65 3.96 1.65 3.96 1.54 4.08 1.54 4.08 1.65 4.845 1.65 4.845 1.54 4.965 1.54 4.965 1.65 6.045 1.65 6.045 1.51 6.105 1.51 6.105 1.65 6.61 1.65 6.61 1.185 6.67 1.185 6.67 1.65 7.55 1.65 7.55 1.345 7.61 1.345 7.61 1.65 8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 0.06 7.555 0.06 7.555 0.555 7.495 0.555 7.495 0.06 6.67 0.06 6.67 0.555 6.61 0.555 6.61 0.06 6.15 0.06 6.15 0.17 6.03 0.17 6.03 0.06 4.965 0.06 4.965 0.55 4.905 0.55 4.905 0.06 2.28 0.06 2.28 0.17 2.16 0.17 2.16 0.06 1.38 0.06 1.38 0.49 1.32 0.49 1.32 0.06 0.555 0.06 0.555 0.635 0.495 0.635 0.495 0.06 0 0.06 0 -0.06 8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.925 1.305 7.865 1.305 7.865 1.245 7.255 1.245 7.255 0.92 7.315 0.92 7.315 1.185 7.865 1.185 7.865 0.525 7.68 0.525 7.68 0.465 7.925 0.465 ;
      POLYGON 7.275 0.55 6.985 0.55 6.985 1.215 7.075 1.215 7.075 1.275 6.925 1.275 6.925 0.715 6.45 0.715 6.45 0.39 5.48 0.39 5.48 0.49 5.605 0.49 5.605 0.755 5.665 0.755 5.665 1.075 5.725 1.075 5.725 1.135 5.605 1.135 5.605 0.815 5.545 0.815 5.545 0.55 5.42 0.55 5.42 0.33 6.51 0.33 6.51 0.655 6.925 0.655 6.925 0.49 7.275 0.49 ;
      POLYGON 6.495 1.245 6.055 1.245 6.055 0.745 5.925 0.745 5.925 0.665 6.055 0.665 6.055 0.49 6.35 0.49 6.35 0.55 6.115 0.55 6.115 1.185 6.495 1.185 ;
      POLYGON 5.94 1.295 4.905 1.295 4.905 1.205 4.51 1.205 4.51 1.075 4.22 1.075 4.22 0.88 4.16 0.88 4.16 0.82 4.28 0.82 4.28 1.015 4.57 1.015 4.57 1.145 4.965 1.145 4.965 1.235 5.445 1.235 5.445 0.975 5.325 0.975 5.325 0.65 5.445 0.65 5.445 0.915 5.505 0.915 5.505 1.235 5.88 1.235 5.88 0.97 5.765 0.97 5.765 0.55 5.705 0.55 5.705 0.49 5.825 0.49 5.825 0.91 5.94 0.91 ;
      POLYGON 5.345 1.135 5.165 1.135 5.165 0.715 4.58 0.715 4.58 0.655 5.165 0.655 5.165 0.49 5.215 0.49 5.215 0.43 5.275 0.43 5.275 0.55 5.225 0.55 5.225 1.075 5.345 1.075 ;
      POLYGON 5.065 0.875 4.73 0.875 4.73 0.985 4.79 0.985 4.79 1.045 4.67 1.045 4.67 0.875 4.42 0.875 4.42 0.68 4.06 0.68 4.06 0.99 3.745 0.99 3.745 0.93 4 0.93 4 0.41 4.06 0.41 4.06 0.62 4.42 0.62 4.42 0.545 4.435 0.545 4.435 0.455 4.495 0.455 4.495 0.59 4.48 0.59 4.48 0.815 5.065 0.815 ;
      POLYGON 4.745 0.55 4.685 0.55 4.685 0.355 4.32 0.355 4.32 0.52 4.2 0.52 4.2 0.46 4.26 0.46 4.26 0.295 4.745 0.295 ;
      POLYGON 4.25 1.395 3.86 1.395 3.86 1.44 2.84 1.44 2.84 1.5 2.78 1.5 2.78 1.44 1.54 1.44 1.54 1.22 1.665 1.22 1.665 0.535 1.64 0.535 1.64 0.395 1.7 0.395 1.7 0.475 1.725 0.475 1.725 1.28 1.6 1.28 1.6 1.38 3.8 1.38 3.8 1.335 4.25 1.335 ;
      POLYGON 4.025 0.31 3.9 0.31 3.9 0.815 3.61 0.815 3.61 0.855 3.53 0.855 3.53 0.735 3.82 0.735 3.82 0.23 4.025 0.23 ;
      POLYGON 3.72 0.635 3.43 0.635 3.43 0.955 3.54 0.955 3.54 1.075 3.48 1.075 3.48 1.015 3.37 1.015 3.37 0.88 2.42 0.88 2.42 0.725 2.15 0.725 2.15 0.785 2.09 0.785 2.09 0.665 2.48 0.665 2.48 0.82 3.37 0.82 3.37 0.575 3.66 0.575 3.66 0.41 3.72 0.41 ;
      POLYGON 3.545 0.475 3.27 0.475 3.27 0.72 2.815 0.72 2.815 0.495 2.875 0.495 2.875 0.66 3.21 0.66 3.21 0.415 3.545 0.415 ;
      RECT 2.505 0.995 3.27 1.075 ;
      POLYGON 3.11 0.56 2.975 0.56 2.975 0.395 2.715 0.395 2.715 0.535 2.7 0.535 2.7 0.56 2.58 0.56 2.58 0.5 2.64 0.5 2.64 0.475 2.655 0.475 2.655 0.335 3.035 0.335 3.035 0.5 3.11 0.5 ;
      POLYGON 2.555 0.375 1.99 0.375 1.99 0.885 2.075 0.885 2.075 1.105 2.015 1.105 2.015 0.945 1.93 0.945 1.93 0.375 1.8 0.375 1.8 0.295 1.54 0.295 1.54 0.65 1.335 0.65 1.335 0.655 1.215 0.655 1.215 0.59 1.48 0.59 1.48 0.235 1.86 0.235 1.86 0.315 2.555 0.315 ;
      POLYGON 0.76 1.02 0.68 1.02 0.68 0.815 0.425 0.815 0.425 0.735 0.68 0.735 0.68 0.54 0.76 0.54 ;
  END
END SDFFNSRXL

MACRO SDFFQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQX1 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.281975 LAYER Metal1 ;
    ANTENNADIFFAREA 2.46425 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.19125 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.9318955 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 94.10196075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.14 1.34 0.08 1.34 0.08 0.73 0.06 0.73 0.06 0.6 0.08 0.6 0.08 0.54 0.14 0.54 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.138889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.165 0.705 3.575 0.705 3.575 0.805 3.55 0.805 3.55 1.005 3.49 1.005 3.49 0.745 3.515 0.745 3.515 0.645 3.685 0.645 3.685 0.585 3.745 0.585 3.745 0.625 4.165 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.21 0.885 3.965 0.885 3.965 1.01 3.835 1.01 3.835 0.805 4.21 0.805 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.23 1.005 3.15 1.005 3.15 0.705 3.035 0.705 3.035 0.625 3.15 0.625 3.15 0.62 3.23 0.62 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.505 1 0.34 1 0.34 1.115 0.26 1.115 0.26 0.92 0.425 0.92 0.425 0.78 0.505 0.78 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.285 1.65 0.285 1.22 0.345 1.22 0.345 1.65 1.085 1.65 1.085 1.49 1.205 1.49 1.205 1.55 1.145 1.55 1.145 1.65 2.1 1.65 2.1 1.51 2.16 1.51 2.16 1.65 3.195 1.65 3.195 1.27 3.255 1.27 3.255 1.65 3.94 1.65 3.94 1.27 4 1.27 4 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 4 0.06 4 0.485 3.94 0.485 3.94 0.06 3.255 0.06 3.255 0.485 3.195 0.485 3.195 0.06 2.17 0.06 2.17 0.17 2.05 0.17 2.05 0.06 1.205 0.06 1.205 0.17 1.085 0.17 1.085 0.06 0.345 0.06 0.345 0.52 0.285 0.52 0.285 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.37 1.17 4.205 1.17 4.205 1.295 4.145 1.295 4.145 1.17 3.675 1.17 3.675 0.805 3.735 0.805 3.735 1.11 4.31 1.11 4.31 0.525 4.145 0.525 4.145 0.39 4.205 0.39 4.205 0.465 4.37 0.465 ;
      POLYGON 3.69 0.485 3.415 0.485 3.415 0.645 3.39 0.645 3.39 1.105 3.415 1.105 3.415 1.27 3.69 1.27 3.69 1.39 3.63 1.39 3.63 1.33 3.355 1.33 3.355 1.165 2.76 1.165 2.76 1.105 2.79 1.105 2.79 0.54 2.85 0.54 2.85 1.105 3.33 1.105 3.33 0.585 3.355 0.585 3.355 0.425 3.63 0.425 3.63 0.365 3.69 0.365 ;
      POLYGON 3.08 1.325 2.6 1.325 2.6 0.83 2.63 0.83 2.63 0.425 1.755 0.425 1.755 0.82 1.695 0.82 1.695 0.365 2.335 0.365 2.335 0.275 2.455 0.275 2.455 0.365 3.05 0.365 3.05 0.485 2.99 0.485 2.99 0.425 2.69 0.425 2.69 0.95 2.66 0.95 2.66 1.265 3.08 1.265 ;
      POLYGON 2.53 0.63 2.5 0.63 2.5 1.16 2.44 1.16 2.44 0.96 2.015 0.96 2.015 0.9 2.44 0.9 2.44 0.63 2.41 0.63 2.41 0.57 2.53 0.57 ;
      POLYGON 2.465 1.385 1.805 1.385 1.805 1.445 1.685 1.445 1.685 1.385 1.315 1.385 1.315 1.29 0.605 1.29 0.605 0.54 0.665 0.54 0.665 1.23 1.315 1.23 1.315 0.78 1.435 0.78 1.435 0.84 1.375 0.84 1.375 1.325 2.465 1.325 ;
      POLYGON 2.295 0.8 1.915 0.8 1.915 1.16 1.855 1.16 1.855 0.57 1.975 0.57 1.975 0.63 1.915 0.63 1.915 0.74 2.295 0.74 ;
      POLYGON 1.71 1.16 1.65 1.16 1.65 1.1 1.535 1.1 1.535 0.44 1.01 0.44 1.01 0.435 0.925 0.435 0.925 0.375 1.045 0.375 1.045 0.38 1.595 0.38 1.595 1.04 1.71 1.04 ;
      POLYGON 1.215 0.79 0.91 0.79 0.91 1.07 0.97 1.07 0.97 1.13 0.85 1.13 0.85 0.595 0.765 0.595 0.765 0.44 0.505 0.44 0.505 0.68 0.3 0.68 0.3 0.82 0.24 0.82 0.24 0.62 0.445 0.62 0.445 0.38 0.825 0.38 0.825 0.535 0.91 0.535 0.91 0.73 1.215 0.73 ;
  END
END SDFFQX1

MACRO SDFFQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQX2 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4798 LAYER Metal1 ;
    ANTENNADIFFAREA 2.72035 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.227475 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.90141775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 86.0995715 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.365 1.29 0.305 1.29 0.305 0.73 0.26 0.73 0.26 0.6 0.305 0.6 0.305 0.37 0.365 0.37 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.861111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.48 0.705 3.835 0.705 3.835 0.845 3.81 0.845 3.81 0.96 3.75 0.96 3.75 0.785 3.775 0.785 3.775 0.645 4.035 0.645 4.035 0.625 4.165 0.625 4.165 0.645 4.48 0.645 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.61 0.975 4.435 0.975 4.435 0.895 4.2 0.895 4.2 0.805 4.61 0.805 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.49 0.92 3.34 0.92 3.34 0.975 3.26 0.975 3.26 0.625 3.34 0.625 3.34 0.79 3.49 0.79 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.61 0.74 1.11 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.1 1.65 0.1 0.9 0.16 0.9 0.16 1.65 0.51 1.65 0.51 1.17 0.57 1.17 0.57 1.65 1.235 1.65 1.235 1.33 1.355 1.33 1.355 1.39 1.295 1.39 1.295 1.65 2.36 1.65 2.36 1.51 2.42 1.51 2.42 1.65 3.455 1.65 3.455 1.235 3.515 1.235 3.515 1.65 4.26 1.65 4.26 1.235 4.32 1.235 4.32 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 4.365 0.06 4.365 0.525 4.305 0.525 4.305 0.06 3.515 0.06 3.515 0.525 3.455 0.525 3.455 0.06 2.45 0.06 2.45 0.17 2.33 0.17 2.33 0.06 1.28 0.06 1.28 0.485 1.34 0.485 1.34 0.545 1.22 0.545 1.22 0.06 0.57 0.06 0.57 0.35 0.51 0.35 0.51 0.06 0.16 0.06 0.16 0.35 0.1 0.35 0.1 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.77 1.135 4.525 1.135 4.525 1.26 4.465 1.26 4.465 1.135 4.04 1.135 4.04 0.94 3.935 0.94 3.935 0.88 4.1 0.88 4.1 1.075 4.71 1.075 4.71 0.545 4.52 0.545 4.52 0.425 4.58 0.425 4.58 0.485 4.77 0.485 ;
      POLYGON 4.055 0.525 3.675 0.525 3.675 0.685 3.65 0.685 3.65 1.075 3.94 1.075 3.94 1.26 3.88 1.26 3.88 1.135 3.14 1.135 3.14 1.155 3.02 1.155 3.02 1.095 3.08 1.095 3.08 0.66 3.05 0.66 3.05 0.54 3.11 0.54 3.11 0.6 3.14 0.6 3.14 1.075 3.59 1.075 3.59 0.625 3.615 0.625 3.615 0.465 3.995 0.465 3.995 0.405 4.055 0.405 ;
      POLYGON 3.34 1.315 2.86 1.315 2.86 0.73 2.89 0.73 2.89 0.44 1.985 0.44 1.985 0.82 1.925 0.82 1.925 0.38 3.31 0.38 3.31 0.525 3.25 0.525 3.25 0.44 2.95 0.44 2.95 0.79 2.92 0.79 2.92 0.89 2.98 0.89 2.98 0.95 2.92 0.95 2.92 1.255 3.34 1.255 ;
      POLYGON 2.79 0.63 2.76 0.63 2.76 1.185 2.7 1.185 2.7 0.975 2.245 0.975 2.245 0.915 2.67 0.915 2.67 0.57 2.79 0.57 ;
      POLYGON 2.725 1.41 2.035 1.41 2.035 1.445 1.915 1.445 1.915 1.41 1.545 1.41 1.545 1.23 0.89 1.23 0.89 1.29 0.83 1.29 0.83 1.17 0.84 1.17 0.84 0.37 0.9 0.37 0.9 1.17 1.545 1.17 1.545 0.805 1.665 0.805 1.665 0.865 1.605 0.865 1.605 1.35 2.725 1.35 ;
      POLYGON 2.545 0.815 2.145 0.815 2.145 1.185 2.085 1.185 2.085 0.57 2.205 0.57 2.205 0.63 2.145 0.63 2.145 0.755 2.545 0.755 ;
      POLYGON 1.94 1.185 1.88 1.185 1.88 1.125 1.765 1.125 1.765 0.705 1.265 0.705 1.265 0.82 1.205 0.82 1.205 0.645 1.765 0.645 1.765 0.54 1.825 0.54 1.825 1.065 1.94 1.065 ;
      POLYGON 1.445 0.98 1.12 0.98 1.12 0.99 1 0.99 1 0.93 1.045 0.93 1.045 0.515 1 0.515 1 0.27 0.74 0.27 0.74 0.51 0.525 0.51 0.525 0.65 0.465 0.65 0.465 0.45 0.68 0.45 0.68 0.21 1.06 0.21 1.06 0.455 1.105 0.455 1.105 0.92 1.445 0.92 ;
  END
END SDFFQX2

MACRO SDFFQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQX4 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.9074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.165 0.705 4.575 0.705 4.575 0.985 4.455 0.985 4.455 0.925 4.515 0.925 4.515 0.645 5.035 0.645 5.035 0.625 5.165 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.205 0.895 4.94 0.895 4.94 1.015 4.835 1.015 4.835 0.805 5.205 0.805 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.355 0.875 4.165 0.875 4.165 0.985 4.085 0.985 4.085 0.895 4.005 0.895 4.005 0.755 4.355 0.755 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.34 0.73 0.31 0.73 0.31 0.97 0.23 0.97 0.23 0.65 0.26 0.65 0.26 0.5 0.34 0.5 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.9456 LAYER Metal1 ;
    ANTENNADIFFAREA 3.23495 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.30915 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.52806075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 75.021834 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.07 0.63 0.935 0.63 0.935 0.885 0.98 0.885 0.98 1.29 0.92 1.29 0.92 0.945 0.875 0.945 0.875 0.66 0.57 0.66 0.57 1.29 0.51 1.29 0.51 0.73 0.46 0.73 0.46 0.6 0.48 0.6 0.48 0.57 0.6 0.57 0.6 0.6 0.875 0.6 0.875 0.57 1.07 0.57 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 1.77 0 1.77 0 1.65 0.305 1.65 0.305 1.07 0.365 1.07 0.365 1.65 0.715 1.65 0.715 0.9 0.775 0.9 0.775 1.65 1.125 1.65 1.125 0.9 1.185 0.9 1.185 1.65 1.565 1.65 1.565 1.155 1.625 1.155 1.625 1.65 2.62 1.65 2.62 1.54 2.74 1.54 2.74 1.65 4.165 1.65 4.165 1.245 4.225 1.245 4.225 1.65 4.91 1.65 4.91 1.275 5.03 1.275 5.03 1.335 4.97 1.335 4.97 1.65 5.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 0.06 5.045 0.06 5.045 0.525 4.985 0.525 4.985 0.06 4.255 0.06 4.255 0.495 4.135 0.495 4.135 0.435 4.195 0.435 4.195 0.06 2.825 0.06 2.825 0.2 2.765 0.2 2.765 0.06 1.75 0.06 1.75 0.2 1.69 0.2 1.69 0.06 1.305 0.06 1.305 0.17 1.185 0.17 1.185 0.06 0.835 0.06 0.835 0.17 0.715 0.17 0.715 0.06 0.335 0.06 0.335 0.2 0.275 0.2 0.275 0.06 0 0.06 0 -0.06 5.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.365 1.175 5.205 1.175 5.205 1.27 5.145 1.27 5.145 1.175 4.675 1.175 4.675 0.99 4.735 0.99 4.735 1.115 5.305 1.115 5.305 0.525 5.2 0.525 5.2 0.405 5.26 0.405 5.26 0.465 5.365 0.465 ;
      POLYGON 4.735 0.545 4.415 0.545 4.415 0.655 3.905 0.655 3.905 1.085 4.575 1.085 4.575 1.27 4.515 1.27 4.515 1.145 3.465 1.145 3.465 1.205 3.405 1.205 3.405 1.085 3.845 1.085 3.845 0.36 3.525 0.36 3.525 0.605 3.405 0.605 3.405 0.545 3.465 0.545 3.465 0.3 3.905 0.3 3.905 0.595 4.355 0.595 4.355 0.485 4.675 0.485 4.675 0.425 4.735 0.425 ;
      POLYGON 4.05 1.335 3.625 1.335 3.625 1.365 3.245 1.365 3.245 1.31 2.225 1.31 2.225 0.925 2.08 0.925 2.08 0.985 2.02 0.985 2.02 0.865 2.285 0.865 2.285 0.805 2.345 0.805 2.345 0.925 2.285 0.925 2.285 1.25 3.245 1.25 3.245 0.895 3.625 0.895 3.625 0.46 3.745 0.46 3.745 0.52 3.685 0.52 3.685 0.955 3.305 0.955 3.305 1.305 3.565 1.305 3.565 1.275 4.05 1.275 ;
      POLYGON 3.46 0.795 3.245 0.795 3.245 0.44 2.985 0.44 2.985 0.96 2.925 0.96 2.925 0.44 1.745 0.44 1.745 0.4 0.13 0.4 0.13 1.02 0.07 1.02 0.07 0.34 1.805 0.34 1.805 0.38 3.305 0.38 3.305 0.735 3.46 0.735 ;
      POLYGON 3.145 1.15 2.765 1.15 2.765 0.98 2.62 0.98 2.62 0.92 2.825 0.92 2.825 1.09 3.085 1.09 3.085 0.54 3.145 0.54 ;
      POLYGON 2.815 0.82 2.755 0.82 2.755 0.76 2.505 0.76 2.505 1.15 2.385 1.15 2.385 1.09 2.445 1.09 2.445 0.54 2.505 0.54 2.505 0.7 2.815 0.7 ;
      POLYGON 2.3 0.63 2.125 0.63 2.125 0.765 1.92 0.765 1.92 1.09 2.1 1.09 2.1 1.15 1.86 1.15 1.86 1.005 1.52 1.005 1.52 0.82 1.58 0.82 1.58 0.945 1.86 0.945 1.86 0.705 2.065 0.705 2.065 0.57 2.3 0.57 ;
      POLYGON 1.76 0.845 1.7 0.845 1.7 0.72 1.42 0.72 1.42 1.29 1.36 1.29 1.36 0.79 1.035 0.79 1.035 0.73 1.36 0.73 1.36 0.5 1.54 0.5 1.54 0.56 1.42 0.56 1.42 0.66 1.76 0.66 ;
  END
END SDFFQX4

MACRO SDFFQXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFQXL 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.42145 LAYER Metal1 ;
    ANTENNADIFFAREA 2.47435 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1782 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.58838375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 104.4444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.41 0.14 1.35 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.4444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.365 0.705 4.235 0.705 4.235 0.685 3.825 0.685 3.825 0.965 3.705 0.965 3.705 0.905 3.765 0.905 3.765 0.625 4.365 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.37 0.94 3.925 0.94 3.925 0.805 4.165 0.805 4.165 0.86 4.37 0.86 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.945 0.815 3.445 0.895 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.41 1.06 0.34 1.06 0.34 1.225 0.26 1.225 0.26 0.98 0.33 0.98 0.33 0.795 0.41 0.795 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.77 0 1.77 0 1.65 0.285 1.65 0.285 1.325 0.345 1.325 0.345 1.65 1.05 1.65 1.05 1.45 1.17 1.45 1.17 1.51 1.11 1.51 1.11 1.65 2.065 1.65 2.065 1.45 2.185 1.45 2.185 1.51 2.125 1.51 2.125 1.65 3.355 1.65 3.355 1.295 3.475 1.295 3.475 1.355 3.415 1.355 3.415 1.65 4.18 1.65 4.18 1.295 4.3 1.295 4.3 1.355 4.24 1.355 4.24 1.65 4.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 0.06 4.27 0.06 4.27 0.525 4.21 0.525 4.21 0.06 3.385 0.06 3.385 0.525 3.325 0.525 3.325 0.06 2.115 0.06 2.115 0.17 1.995 0.17 1.995 0.06 1.17 0.06 1.17 0.17 1.05 0.17 1.05 0.06 0.305 0.06 0.305 0.2 0.245 0.2 0.245 0.06 0 0.06 0 -0.06 4.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.53 1.29 4.415 1.29 4.415 1.1 3.925 1.1 3.925 1.04 4.47 1.04 4.47 0.43 4.53 0.43 ;
      POLYGON 3.96 0.525 3.665 0.525 3.665 0.78 3.605 0.78 3.605 1.065 3.825 1.065 3.825 1.2 3.86 1.2 3.86 1.32 3.8 1.32 3.8 1.26 3.765 1.26 3.765 1.125 2.785 1.125 2.785 0.57 2.905 0.57 2.905 0.63 2.845 0.63 2.845 1.065 3.545 1.065 3.545 0.72 3.605 0.72 3.605 0.465 3.9 0.465 3.9 0.405 3.96 0.405 ;
      POLYGON 3.255 1.285 2.625 1.285 2.625 0.445 1.72 0.445 1.72 0.82 1.66 0.82 1.66 0.385 2.34 0.385 2.34 0.25 2.46 0.25 2.46 0.385 3.15 0.385 3.15 0.435 3.21 0.435 3.21 0.495 3.09 0.495 3.09 0.445 2.685 0.445 2.685 1.225 3.255 1.225 ;
      POLYGON 2.525 0.63 2.465 0.63 2.465 0.93 2.525 0.93 2.525 1.125 2.465 1.125 2.465 0.99 2.04 0.99 2.04 0.925 1.98 0.925 1.98 0.865 2.1 0.865 2.1 0.93 2.405 0.93 2.405 0.57 2.525 0.57 ;
      POLYGON 2.49 1.35 1.74 1.35 1.74 1.445 1.62 1.445 1.62 1.35 0.51 1.35 0.51 0.465 0.63 0.465 0.63 0.525 0.57 0.525 0.57 1.29 1.28 1.29 1.28 0.745 1.4 0.745 1.4 0.805 1.34 0.805 1.34 1.29 2.49 1.29 ;
      POLYGON 2.26 0.83 2.2 0.83 2.2 0.765 1.88 0.765 1.88 1.095 1.76 1.095 1.76 1.035 1.82 1.035 1.82 0.545 1.94 0.545 1.94 0.605 1.88 0.605 1.88 0.705 2.26 0.705 ;
      POLYGON 1.645 1.125 1.585 1.125 1.585 0.98 1.5 0.98 1.5 0.435 0.89 0.435 0.89 0.375 1.56 0.375 1.56 0.92 1.645 0.92 ;
      POLYGON 1.18 0.79 0.875 0.79 0.875 1.035 0.935 1.035 0.935 1.095 0.815 1.095 0.815 0.595 0.73 0.595 0.73 0.365 0.41 0.365 0.41 0.695 0.24 0.695 0.24 0.635 0.35 0.635 0.35 0.305 0.79 0.305 0.79 0.535 0.875 0.535 0.875 0.73 1.18 0.73 ;
  END
END SDFFQXL

MACRO SDFFRHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRHQX1 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.83605 LAYER Metal1 ;
    ANTENNADIFFAREA 3.109175 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2601 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.903691 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 87.5432525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.175 1.41 0.115 1.41 0.115 0.73 0.06 0.73 0.06 0.6 0.115 0.6 0.115 0.31 0.175 0.31 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.55775575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.63 0.765 4.57 0.765 4.57 0.705 3.98 0.705 3.98 1 3.92 1 3.92 0.625 4.585 0.625 4.585 0.645 4.63 0.645 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.87179475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.26 0.79 4.48 1.045 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.79487175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.65 0.645 3.74 0.925 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.750809 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.17 0.77 1.37 0.995 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.4074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.235 0.815 0.5 0.95 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.32 1.65 0.32 1.05 0.38 1.05 0.38 1.65 0.745 1.65 0.745 1.395 0.865 1.395 0.865 1.475 0.805 1.475 0.805 1.65 1.275 1.65 1.275 1.235 1.335 1.235 1.335 1.65 2.22 1.65 2.22 1.475 2.16 1.475 2.16 1.395 2.28 1.395 2.28 1.65 2.63 1.65 2.63 1.52 2.75 1.52 2.75 1.65 3.59 1.65 3.59 1.49 3.65 1.49 3.65 1.65 4.335 1.65 4.335 1.3 4.395 1.3 4.395 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 4.5 0.06 4.5 0.525 4.44 0.525 4.44 0.06 3.68 0.06 3.68 0.565 3.62 0.565 3.62 0.06 2.28 0.06 2.28 0.435 2.22 0.435 2.22 0.06 1.275 0.06 1.275 0.23 1.335 0.23 1.335 0.29 1.215 0.29 1.215 0.06 0.38 0.06 0.38 0.55 0.32 0.55 0.32 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.75 1.205 4.705 1.205 4.705 1.265 4.645 1.265 4.645 1.205 4.09 1.205 4.09 0.89 4.15 0.89 4.15 1.145 4.69 1.145 4.69 0.55 4.645 0.55 4.645 0.43 4.705 0.43 4.705 0.49 4.75 0.49 ;
      POLYGON 4.19 0.545 3.86 0.545 3.86 1.1 3.99 1.1 3.99 1.44 3.93 1.44 3.93 1.3 3.215 1.3 3.215 0.81 2.995 0.81 2.995 0.42 3.115 0.42 3.115 0.48 3.055 0.48 3.055 0.75 3.275 0.75 3.275 1.24 3.8 1.24 3.8 0.485 4.13 0.485 4.13 0.425 4.19 0.425 ;
      POLYGON 3.52 1.44 2.635 1.44 2.635 1.33 1.52 1.33 1.52 1.155 1.215 1.155 1.215 1.315 0.56 1.315 0.56 0.45 0.62 0.45 0.62 1.255 1.155 1.255 1.155 1.095 1.52 1.095 1.52 0.67 1.58 0.67 1.58 1.27 1.82 1.27 1.82 0.875 1.88 0.875 1.88 1.27 2.695 1.27 2.695 1.38 3.52 1.38 ;
      POLYGON 3.475 1.18 3.415 1.18 3.415 0.65 3.155 0.65 3.155 0.59 3.215 0.59 3.215 0.32 2.715 0.32 2.715 0.595 2.735 0.595 2.735 0.715 2.655 0.715 2.655 0.585 2.1 0.585 2.1 0.31 1.88 0.31 1.88 0.675 1.82 0.675 1.82 0.25 2.16 0.25 2.16 0.525 2.655 0.525 2.655 0.26 3.275 0.26 3.275 0.59 3.415 0.59 3.415 0.455 3.475 0.455 ;
      POLYGON 3.07 1.21 3.01 1.21 3.01 0.97 2.09 0.97 2.09 0.84 2.15 0.84 2.15 0.91 2.835 0.91 2.835 0.48 2.775 0.48 2.775 0.42 2.895 0.42 2.895 0.91 3.07 0.91 ;
      RECT 2.395 1.1 2.895 1.16 ;
      POLYGON 2.555 0.8 2.495 0.8 2.495 0.705 2.005 0.705 2.005 1.185 1.945 1.185 1.945 0.39 2.005 0.39 2.005 0.645 2.555 0.645 ;
      POLYGON 1.74 1.185 1.68 1.185 1.68 0.45 0.94 0.45 0.94 0.68 0.88 0.68 0.88 0.39 1.68 0.39 1.68 0.33 1.74 0.33 ;
      POLYGON 1.4 0.67 1.07 0.67 1.07 1.185 1.01 1.185 1.01 0.84 0.76 0.84 0.76 0.35 0.5 0.35 0.5 0.69 0.335 0.69 0.335 0.75 0.275 0.75 0.275 0.63 0.44 0.63 0.44 0.29 0.82 0.29 0.82 0.78 1.01 0.78 1.01 0.61 1.34 0.61 1.34 0.55 1.4 0.55 ;
  END
END SDFFRHQX1

MACRO SDFFRHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRHQX2 0 0 ;
  SIZE 5.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1616 LAYER Metal1 ;
    ANTENNADIFFAREA 3.74445 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.28935 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.9265595 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 84.98704 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.34 1.315 0.26 1.315 0.26 1.005 0.255 1.005 0.255 0.42 0.335 0.42 0.335 0.925 0.34 0.925 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.56765675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.475 0.715 5.14 0.715 5.14 0.705 4.84 0.705 4.84 0.915 4.78 0.915 4.78 0.645 5.035 0.645 5.035 0.625 5.165 0.625 5.165 0.645 5.2 0.645 5.2 0.655 5.475 0.655 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.61 0.925 5.14 0.925 5.14 0.845 5.195 0.845 5.195 0.815 5.61 0.815 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.52 0.87 4.44 0.87 4.44 0.68 4.34 0.68 4.34 0.73 4.26 0.73 4.26 0.6 4.52 0.6 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.75404525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.855 0.995 1.48 0.995 1.48 0.79 1.665 0.79 1.665 0.815 1.855 0.815 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 1.095 0.66 1.095 0.66 0.92 0.595 0.92 0.595 0.66 0.74 0.66 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 1.77 0 1.77 0 1.65 0.075 1.65 0.075 0.925 0.135 0.925 0.135 1.65 0.485 1.65 0.485 1.195 0.545 1.195 0.545 1.65 1.265 1.65 1.265 1.415 1.325 1.415 1.325 1.65 1.765 1.65 1.765 1.475 1.705 1.475 1.705 1.415 1.825 1.415 1.825 1.65 2.89 1.65 2.89 1.475 2.83 1.475 2.83 1.415 2.95 1.415 2.95 1.65 3.3 1.65 3.3 1.54 3.42 1.54 3.42 1.65 4.4 1.65 4.4 1.54 4.52 1.54 4.52 1.65 5.225 1.65 5.225 1.235 5.285 1.235 5.285 1.65 5.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 0.06 5.36 0.06 5.36 0.545 5.3 0.545 5.3 0.06 4.52 0.06 4.52 0.435 4.46 0.435 4.46 0.06 3.095 0.06 3.095 0.17 2.975 0.17 2.975 0.06 1.71 0.06 1.71 0.25 1.77 0.25 1.77 0.31 1.65 0.31 1.65 0.06 0.54 0.06 0.54 0.4 0.48 0.4 0.48 0.06 0.13 0.06 0.13 0.4 0.07 0.4 0.07 0.06 0 0.06 0 -0.06 5.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.77 1.085 5.52 1.085 5.52 1.145 5.46 1.145 5.46 1.085 4.98 1.085 4.98 0.805 5.04 0.805 5.04 1.025 5.71 1.025 5.71 0.555 5.515 0.555 5.515 0.435 5.575 0.435 5.575 0.495 5.77 0.495 ;
      POLYGON 4.965 0.545 4.68 0.545 4.68 1.015 4.88 1.015 4.88 1.355 4.82 1.355 4.82 1.075 4.475 1.075 4.475 1.215 3.94 1.215 3.94 0.875 3.82 0.875 3.82 0.44 3.94 0.44 3.94 0.5 3.88 0.5 3.88 0.815 4 0.815 4 1.155 4.415 1.155 4.415 1.015 4.62 1.015 4.62 0.485 4.905 0.485 4.905 0.425 4.965 0.425 ;
      POLYGON 4.36 1.375 3.33 1.375 3.33 1.335 3.05 1.335 3.05 1.315 0.69 1.315 0.69 1.195 0.84 1.195 0.84 0.57 0.8 0.57 0.8 0.42 0.86 0.42 0.86 0.51 0.9 0.51 0.9 1.255 1.955 1.255 1.955 0.69 2.015 0.69 2.015 1.255 2.275 1.255 2.275 0.82 2.335 0.82 2.335 1.255 3.11 1.255 3.11 1.275 3.39 1.275 3.39 1.315 4.36 1.315 ;
      POLYGON 4.315 1.055 4.1 1.055 4.1 0.715 3.98 0.715 3.98 0.655 4.1 0.655 4.1 0.34 3.5 0.34 3.5 0.6 3.52 0.6 3.52 0.72 3.44 0.72 3.44 0.34 2.495 0.34 2.495 0.6 2.555 0.6 2.555 0.66 2.435 0.66 2.435 0.28 4.16 0.28 4.16 0.995 4.315 0.995 ;
      POLYGON 3.795 1.215 3.735 1.215 3.735 1.035 3.66 1.035 3.66 0.88 3.12 0.88 3.12 0.78 2.815 0.78 2.815 0.72 3.18 0.72 3.18 0.82 3.66 0.82 3.66 0.5 3.6 0.5 3.6 0.44 3.72 0.44 3.72 0.975 3.795 0.975 ;
      POLYGON 3.57 1.215 3.49 1.215 3.49 1.175 3.21 1.175 3.21 1.155 3.065 1.155 3.065 1.075 3.29 1.075 3.29 1.095 3.57 1.095 ;
      POLYGON 3.34 0.69 3.28 0.69 3.28 0.62 2.715 0.62 2.715 1.07 2.595 1.07 2.595 1.01 2.655 1.01 2.655 0.5 2.595 0.5 2.595 0.44 2.715 0.44 2.715 0.56 3.34 0.56 ;
      POLYGON 2.175 1.155 2.115 1.155 2.115 0.47 1.22 0.47 1.22 0.7 1.16 0.7 1.16 0.41 2.115 0.41 2.115 0.35 2.175 0.35 ;
      POLYGON 1.835 0.69 1.38 0.69 1.38 1.095 1.59 1.095 1.59 1.155 1.32 1.155 1.32 0.86 1 0.86 1 0.32 0.7 0.32 0.7 0.56 0.495 0.56 0.495 0.71 0.435 0.71 0.435 0.5 0.64 0.5 0.64 0.26 1.06 0.26 1.06 0.8 1.32 0.8 1.32 0.63 1.775 0.63 1.775 0.57 1.835 0.57 ;
  END
END SDFFRHQX2

MACRO SDFFRHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRHQX4 0 0 ;
  SIZE 7.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.29372925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.965 0.705 6.835 0.705 6.835 0.555 6.3 0.555 6.3 0.665 6.18 0.665 6.18 0.495 6.895 0.495 6.895 0.625 6.965 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.735 0.96 6.46 0.96 6.46 0.79 6.655 0.79 6.655 0.655 6.735 0.655 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.895 0.88 5.815 0.88 5.815 0.705 5.57 0.705 5.57 0.625 5.895 0.625 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.069525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 15.6850055 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.93 0.905 3.54 0.905 3.54 0.395 2.265 0.395 2.265 0.745 2.205 0.745 2.205 0.395 1.775 0.395 1.775 0.755 1.66 0.755 1.66 0.6 1.715 0.6 1.715 0.335 3.6 0.335 3.6 0.845 3.87 0.845 3.87 0.76 3.93 0.76 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.685 0.34 1.185 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.723 LAYER Metal1 ;
    ANTENNADIFFAREA 4.9105 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.371025 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.03436425 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 77.533859 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.36 0.61 1.285 0.61 1.285 1.02 1.165 1.02 1.165 0.96 1.225 0.96 1.225 0.66 0.94 0.66 0.94 1.02 0.695 1.02 0.695 0.96 0.88 0.96 0.88 0.73 0.86 0.73 0.86 0.52 0.94 0.52 0.94 0.6 1.225 0.6 1.225 0.55 1.36 0.55 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 1.77 0 1.77 0 1.65 0.46 1.65 0.46 1.455 0.58 1.455 0.58 1.515 0.52 1.515 0.52 1.65 0.93 1.65 0.93 1.455 1.05 1.455 1.05 1.515 0.99 1.515 0.99 1.65 1.45 1.65 1.45 1.455 1.57 1.455 1.57 1.515 1.51 1.515 1.51 1.65 1.95 1.65 1.95 1.51 2.01 1.51 2.01 1.65 2.42 1.65 2.42 1.51 2.48 1.51 2.48 1.65 3.735 1.65 3.735 1.54 3.855 1.54 3.855 1.65 4.425 1.65 4.425 1.54 4.545 1.54 4.545 1.65 5.79 1.65 5.79 1.165 5.85 1.165 5.85 1.65 6.515 1.65 6.515 1.22 6.575 1.22 6.575 1.65 7.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 0.06 6.575 0.06 6.575 0.395 6.515 0.395 6.515 0.06 5.79 0.06 5.79 0.305 5.85 0.305 5.85 0.365 5.73 0.365 5.73 0.06 3.795 0.06 3.795 0.5 3.735 0.5 3.735 0.06 2.51 0.06 2.51 0.17 2.39 0.17 2.39 0.06 1.615 0.06 1.615 0.5 1.555 0.5 1.555 0.06 1.125 0.06 1.125 0.5 1.065 0.5 1.065 0.06 0.715 0.06 0.715 0.5 0.655 0.5 0.655 0.06 0 0.06 0 -0.06 7.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.125 1.12 6.3 1.12 6.3 0.88 5.995 0.88 5.995 0.65 6.055 0.65 6.055 0.82 6.36 0.82 6.36 1.06 7.065 1.06 7.065 0.525 6.995 0.525 6.995 0.405 7.055 0.405 7.055 0.465 7.125 0.465 ;
      POLYGON 6.2 1.34 6.14 1.34 6.14 1.04 5.41 1.04 5.41 1.025 5.285 1.025 5.285 0.965 5.41 0.965 5.41 0.345 4.91 0.345 4.91 0.5 4.85 0.5 4.85 0.285 5.47 0.285 5.47 0.465 5.95 0.465 5.95 0.335 6.16 0.335 6.16 0.395 6.01 0.395 6.01 0.525 5.47 0.525 5.47 0.98 6.2 0.98 ;
      POLYGON 5.69 1.445 4.645 1.445 4.645 1.385 1.67 1.385 1.67 1.355 0.1 1.355 0.1 0.525 0.4 0.525 0.4 0.585 0.16 0.585 0.16 1.295 1.73 1.295 1.73 1.325 4.705 1.325 4.705 1.385 5.69 1.385 ;
      POLYGON 5.585 1.26 4.805 1.26 4.805 1.225 3.16 1.225 3.16 0.89 2.905 0.89 2.905 0.77 2.965 0.77 2.965 0.83 3.16 0.83 3.16 0.69 3.28 0.69 3.28 0.75 3.22 0.75 3.22 1.165 4.805 1.165 4.805 0.835 4.55 0.835 4.55 0.775 4.865 0.775 4.865 1.2 5.125 1.2 5.125 0.445 5.31 0.445 5.31 0.505 5.185 0.505 5.185 1.2 5.525 1.2 5.525 1.14 5.585 1.14 ;
      POLYGON 5.025 1.055 4.965 1.055 4.965 0.66 3.76 0.66 3.76 0.745 3.7 0.745 3.7 0.6 4.645 0.6 4.645 0.465 4.705 0.465 4.705 0.6 5.025 0.6 ;
      POLYGON 4.705 1.055 4.19 1.055 4.19 0.975 4.625 0.975 4.625 0.935 4.705 0.935 ;
      POLYGON 4.375 0.86 4.09 0.86 4.09 1.065 3.32 1.065 3.32 1.005 3.38 1.005 3.38 0.555 3.32 0.555 3.32 0.495 3.44 0.495 3.44 1.005 4.03 1.005 4.03 0.8 4.375 0.8 ;
      POLYGON 3.215 0.555 3.06 0.555 3.06 0.67 2.805 0.67 2.805 0.99 3.015 0.99 3.015 1.225 2.955 1.225 2.955 1.05 2.745 1.05 2.745 0.67 2.425 0.67 2.425 0.905 2.035 0.905 2.035 0.735 2.095 0.735 2.095 0.845 2.365 0.845 2.365 0.61 3 0.61 3 0.495 3.215 0.495 ;
      POLYGON 2.645 0.86 2.585 0.86 2.585 1.065 2.245 1.065 2.245 1.125 2.185 1.125 2.185 1.065 1.445 1.065 1.445 0.86 1.385 0.86 1.385 0.8 1.505 0.8 1.505 1.005 1.875 1.005 1.875 0.495 2.01 0.495 2.01 0.555 1.935 0.555 1.935 1.005 2.525 1.005 2.525 0.8 2.645 0.8 ;
  END
END SDFFRHQX4

MACRO SDFFRHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRHQX8 0 0 ;
  SIZE 7.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.16171625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.565 0.715 7.345 0.715 7.345 0.705 6.84 0.705 6.84 0.915 6.78 0.915 6.78 0.645 7.345 0.645 7.345 0.625 7.565 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.61 0.895 7.365 0.895 7.365 0.915 7.13 0.915 7.13 0.815 7.61 0.815 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.52 0.895 6.44 0.895 6.44 0.705 6.34 0.705 6.34 0.73 6.26 0.73 6.26 0.6 6.34 0.6 6.34 0.625 6.52 0.625 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.655 0.915 3.4 0.915 3.4 0.815 3.545 0.815 3.545 0.59 3.655 0.59 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1161 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.110925 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.04665325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.8749155 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.545 0.755 2.39 0.755 2.39 0.405 1.965 0.405 1.965 0.765 1.805 0.765 1.805 0.705 1.835 0.705 1.835 0.625 1.905 0.625 1.905 0.345 2.45 0.345 2.45 0.695 2.545 0.695 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3068 LAYER Metal1 ;
    ANTENNADIFFAREA 5.327475 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.528525 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.14871575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 63.8285795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.57 0.66 1.485 0.66 1.485 1.35 1.425 1.35 1.425 0.73 1.075 0.73 1.075 1.35 1.015 1.35 1.015 0.73 0.665 0.73 0.665 1.35 0.605 1.35 0.605 0.73 0.255 0.73 0.255 1.35 0.195 1.35 0.195 0.67 0.26 0.67 0.26 0.54 0.34 0.54 0.34 0.67 0.69 0.67 0.69 0.54 0.75 0.54 0.75 0.67 1.1 0.67 1.1 0.54 1.16 0.54 1.16 0.67 1.425 0.67 1.425 0.6 1.51 0.6 1.51 0.54 1.57 0.54 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.8 1.77 0 1.77 0 1.65 0.4 1.65 0.4 0.905 0.46 0.905 0.46 1.65 0.81 1.65 0.81 0.905 0.87 0.905 0.87 1.65 1.22 1.65 1.22 0.905 1.28 0.905 1.28 1.65 1.66 1.65 1.66 1.175 1.72 1.175 1.72 1.65 2.07 1.65 2.07 1.175 2.13 1.175 2.13 1.65 2.5 1.65 2.5 1.235 2.52 1.235 2.52 1.175 2.58 1.175 2.58 1.295 2.56 1.295 2.56 1.65 2.96 1.65 2.96 1.54 3.08 1.54 3.08 1.65 3.535 1.65 3.535 1.54 3.655 1.54 3.655 1.65 4.715 1.65 4.715 1.135 4.775 1.135 4.775 1.65 5.24 1.65 5.24 1.54 5.36 1.54 5.36 1.65 6.4 1.65 6.4 1.54 6.52 1.54 6.52 1.65 7.215 1.65 7.215 1.235 7.275 1.235 7.275 1.65 7.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.8 0.06 7.36 0.06 7.36 0.525 7.3 0.525 7.3 0.06 6.52 0.06 6.52 0.435 6.46 0.435 6.46 0.06 4.895 0.06 4.895 0.335 4.775 0.335 4.775 0.275 4.835 0.275 4.835 0.06 3.74 0.06 3.74 0.17 3.62 0.17 3.62 0.06 2.61 0.06 2.61 0.485 2.55 0.485 2.55 0.06 1.775 0.06 1.775 0.485 1.715 0.485 1.715 0.06 1.365 0.06 1.365 0.485 1.305 0.485 1.305 0.06 0.955 0.06 0.955 0.485 0.895 0.485 0.895 0.06 0.545 0.06 0.545 0.485 0.485 0.485 0.485 0.06 0 0.06 0 -0.06 7.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.77 1.075 7.51 1.075 7.51 1.135 7.45 1.135 7.45 1.075 6.97 1.075 6.97 0.805 7.03 0.805 7.03 1.015 7.71 1.015 7.71 0.525 7.615 0.525 7.615 0.405 7.675 0.405 7.675 0.465 7.77 0.465 ;
      POLYGON 7.05 0.545 6.68 0.545 6.68 1.015 6.87 1.015 6.87 1.355 6.81 1.355 6.81 1.075 6.445 1.075 6.445 1.215 5.94 1.215 5.94 0.845 5.705 0.845 5.705 0.455 5.825 0.455 5.825 0.515 5.765 0.515 5.765 0.785 6 0.785 6 1.155 6.385 1.155 6.385 1.015 6.62 1.015 6.62 0.485 6.99 0.485 6.99 0.425 7.05 0.425 ;
      POLYGON 6.36 1.385 4.875 1.385 4.875 1.035 4.615 1.035 4.615 1.225 3.915 1.225 3.915 0.49 3.3 0.49 3.3 1.015 3.56 1.015 3.56 1.075 3.24 1.075 3.24 0.43 3.975 0.43 3.975 1.165 4.235 1.165 4.235 0.775 4.295 0.775 4.295 1.165 4.555 1.165 4.555 0.975 4.935 0.975 4.935 1.325 6.36 1.325 ;
      POLYGON 6.285 1.055 6.1 1.055 6.1 0.685 5.865 0.685 5.865 0.625 5.925 0.625 5.925 0.335 5.385 0.335 5.385 0.595 5.395 0.595 5.395 0.715 5.325 0.715 5.325 0.495 4.615 0.495 4.615 0.355 4.295 0.355 4.295 0.615 4.355 0.615 4.355 0.675 4.235 0.675 4.235 0.295 4.675 0.295 4.675 0.435 5.325 0.435 5.325 0.275 5.985 0.275 5.985 0.625 6.1 0.625 6.1 0.455 6.16 0.455 6.16 0.995 6.285 0.995 ;
      POLYGON 5.795 1.225 5.735 1.225 5.735 1.005 5.545 1.005 5.545 0.875 5.005 0.875 5.005 0.84 4.615 0.84 4.615 0.78 5.065 0.78 5.065 0.815 5.545 0.815 5.545 0.495 5.485 0.495 5.485 0.435 5.605 0.435 5.605 0.945 5.795 0.945 ;
      POLYGON 5.59 1.225 5.035 1.225 5.035 1.105 5.115 1.105 5.115 1.145 5.51 1.145 5.51 1.105 5.59 1.105 ;
      POLYGON 5.225 0.715 5.165 0.715 5.165 0.655 4.515 0.655 4.515 0.835 4.455 0.835 4.455 1.065 4.395 1.065 4.395 0.775 4.455 0.775 4.455 0.515 4.395 0.515 4.395 0.455 4.515 0.455 4.515 0.595 5.225 0.595 ;
      POLYGON 4.56 1.46 3.755 1.46 3.755 1.425 2.66 1.425 2.66 1.365 3.815 1.365 3.815 1.4 4.56 1.4 ;
      POLYGON 4.135 1.065 4.075 1.065 4.075 0.33 2.77 0.33 2.77 0.695 2.91 0.695 2.91 0.755 2.77 0.755 2.77 0.915 2.23 0.915 2.23 0.735 2.29 0.735 2.29 0.855 2.71 0.855 2.71 0.27 4.135 0.27 ;
      POLYGON 3.815 1.235 3.01 1.235 3.01 1.075 2.815 1.075 2.815 1.135 2.755 1.135 2.755 1.075 2.365 1.075 2.365 1.295 2.305 1.295 2.305 1.075 1.925 1.075 1.925 1.295 1.865 1.295 1.865 0.965 1.645 0.965 1.645 0.835 1.585 0.835 1.585 0.775 1.705 0.775 1.705 0.905 1.925 0.905 1.925 1.015 2.07 1.015 2.07 0.505 2.13 0.505 2.13 1.015 3.01 1.015 3.01 0.595 2.87 0.595 2.87 0.535 3.07 0.535 3.07 1.175 3.755 1.175 3.755 0.75 3.815 0.75 ;
  END
END SDFFRHQX8

MACRO SDFFRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRX1 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3264 LAYER Metal1 ;
    ANTENNADIFFAREA 3.664625 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2367 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.053232 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 107.07224325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 1.33 0.88 1.33 0.88 0.73 0.86 0.73 0.86 0.6 0.865 0.6 0.865 0.54 0.94 0.54 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3264 LAYER Metal1 ;
    ANTENNADIFFAREA 3.664625 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2367 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.053232 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 107.07224325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.29 1.29 0.21 1.29 0.21 0.73 0.06 0.73 0.06 0.6 0.21 0.6 0.21 0.54 0.29 0.54 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.212963 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.14 0.73 6.06 0.73 6.06 0.525 5.465 0.525 5.465 0.735 5.2 0.735 5.2 0.795 5.14 0.795 5.14 0.675 5.405 0.675 5.405 0.465 6.12 0.465 6.12 0.6 6.14 0.6 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.96 0.745 5.645 0.745 5.645 0.81 5.565 0.81 5.565 0.625 5.96 0.625 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.88 0.575 4.74 0.575 4.74 0.855 4.66 0.855 4.66 0.495 4.88 0.495 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0912 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.81481475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 34.62962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.155 0.815 1.965 0.815 1.965 0.96 1.8 0.96 1.8 0.735 2.155 0.735 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.28 1.11 1.06 1.11 1.06 0.98 1.2 0.98 1.2 0.75 1.28 0.75 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 1.77 0 1.77 0 1.65 0.465 1.65 0.465 1.285 0.525 1.285 0.525 1.65 1.085 1.65 1.085 1.21 1.145 1.21 1.145 1.65 1.75 1.65 1.75 1.51 1.81 1.51 1.81 1.65 2.12 1.65 2.12 1.54 2.24 1.54 2.24 1.65 3.2 1.65 3.2 1.54 3.32 1.54 3.32 1.65 3.67 1.65 3.67 1.38 3.79 1.38 3.79 1.44 3.73 1.44 3.73 1.65 4.795 1.65 4.795 1.51 4.855 1.51 4.855 1.65 5.64 1.65 5.64 1.07 5.7 1.07 5.7 1.65 6.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 0.06 5.67 0.06 5.67 0.305 5.73 0.305 5.73 0.365 5.61 0.365 5.61 0.06 4.785 0.06 4.785 0.395 4.725 0.395 4.725 0.06 3.42 0.06 3.42 0.25 3.3 0.25 3.3 0.19 3.36 0.19 3.36 0.06 2.21 0.06 2.21 0.315 2.15 0.315 2.15 0.06 1.1 0.06 1.1 0.43 1.16 0.43 1.16 0.49 1.04 0.49 1.04 0.06 0.525 0.06 0.525 0.2 0.465 0.2 0.465 0.06 0 0.06 0 -0.06 6.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.3 0.97 6.195 0.97 6.195 1.095 6.135 1.095 6.135 0.97 5.365 0.97 5.365 0.905 5.305 0.905 5.305 0.845 5.425 0.845 5.425 0.91 6.24 0.91 6.24 0.5 6.22 0.5 6.22 0.3 6.28 0.3 6.28 0.44 6.3 0.44 ;
      POLYGON 5.42 0.365 5.04 0.365 5.04 1.07 5.36 1.07 5.36 1.13 5.04 1.13 5.04 1.225 4.24 1.225 4.24 0.93 4.18 0.93 4.18 0.5 4.055 0.5 4.055 0.38 4.115 0.38 4.115 0.44 4.24 0.44 4.24 0.87 4.3 0.87 4.3 1.165 4.98 1.165 4.98 0.305 5.42 0.305 ;
      POLYGON 4.695 1.385 4.08 1.385 4.08 1.28 3.98 1.28 3.98 1.34 3.92 1.34 3.92 1.28 1.38 1.28 1.38 0.97 1.42 0.97 1.42 0.57 1.54 0.57 1.54 0.63 1.48 0.63 1.48 1.03 1.44 1.03 1.44 1.22 2.425 1.22 2.425 0.645 2.485 0.645 2.485 1.22 2.805 1.22 2.805 0.865 2.745 0.865 2.745 0.805 2.865 0.805 2.865 1.22 4.14 1.22 4.14 1.325 4.695 1.325 ;
      POLYGON 4.62 1.065 4.5 1.065 4.5 0.44 4.4 0.44 4.4 0.77 4.34 0.77 4.34 0.28 3.58 0.28 3.58 0.41 3.14 0.41 3.14 0.28 2.805 0.28 2.805 0.66 2.745 0.66 2.745 0.22 3.2 0.22 3.2 0.35 3.52 0.35 3.52 0.22 4.4 0.22 4.4 0.38 4.56 0.38 4.56 1.005 4.62 1.005 ;
      POLYGON 4.095 1.115 4.035 1.115 4.035 1.04 4.02 1.04 4.02 0.85 3.185 0.85 3.185 0.73 3.245 0.73 3.245 0.79 3.85 0.79 3.85 0.38 3.91 0.38 3.91 0.79 4.08 0.79 4.08 0.995 4.095 0.995 ;
      RECT 3.42 0.95 3.92 1.03 ;
      POLYGON 3.695 0.63 3.085 0.63 3.085 1.025 2.965 1.025 2.965 0.965 2.98 0.965 2.98 0.38 3.04 0.38 3.04 0.57 3.695 0.57 ;
      RECT 1.96 1.38 3.48 1.44 ;
      POLYGON 2.705 1.025 2.585 1.025 2.585 0.475 1.86 0.475 1.86 0.28 1.8 0.28 1.8 0.22 1.92 0.22 1.92 0.415 2.585 0.415 2.585 0.355 2.645 0.355 2.645 0.965 2.705 0.965 ;
      POLYGON 2.315 0.695 2.255 0.695 2.255 0.635 1.7 0.635 1.7 1.06 2.005 1.06 2.005 1.12 1.64 1.12 1.64 0.44 1.32 0.44 1.32 0.65 1.1 0.65 1.1 0.82 1.04 0.82 1.04 0.59 1.26 0.59 1.26 0.38 1.71 0.38 1.71 0.575 2.315 0.575 ;
      POLYGON 0.725 1.02 0.645 1.02 0.645 0.81 0.39 0.81 0.39 0.73 0.645 0.73 0.645 0.54 0.725 0.54 ;
  END
END SDFFRX1

MACRO SDFFRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRX2 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.3013 LAYER Metal1 ;
    ANTENNADIFFAREA 3.8091 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.302175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.92512625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 84.43286175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.175 0.99 1.055 0.99 1.055 0.49 1.135 0.49 1.135 0.6 1.14 0.6 1.14 0.73 1.135 0.73 1.135 0.91 1.175 0.91 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.34515 LAYER Metal1 ;
    ANTENNADIFFAREA 3.8091 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.302175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.07024075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 85.053363 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 0.73 0.73 0.73 0.73 0.99 0.56 0.99 0.56 0.91 0.65 0.91 0.65 0.49 0.73 0.49 0.73 0.6 0.74 0.6 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.7314815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.14 0.73 6.06 0.73 6.06 0.68 5.715 0.68 5.715 0.88 5.635 0.88 5.635 0.6 6.14 0.6 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.935 0.86 5.895 0.86 5.895 1.085 5.635 1.085 5.635 1.005 5.815 1.005 5.815 0.78 5.935 0.78 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.215 0.87 5.14 0.87 5.14 1.025 5.06 1.025 5.06 0.79 5.135 0.79 5.135 0.6 5.215 0.6 ;
    END
  END SI
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.039375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 15.1238095 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.77 1.44 2.78 1.44 2.78 1.11 2.46 1.11 2.46 0.9 2.385 0.9 2.385 0.84 2.52 0.84 2.52 0.98 2.54 0.98 2.54 1.05 2.84 1.05 2.84 1.38 3.77 1.38 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.64 0.705 1.515 0.705 1.515 0.945 1.435 0.945 1.435 0.57 1.64 0.57 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 1.77 0 1.77 0 1.65 0.3 1.65 0.3 1.25 0.42 1.25 0.42 1.31 0.36 1.31 0.36 1.65 0.795 1.65 0.795 1.25 0.915 1.25 0.915 1.31 0.855 1.31 0.855 1.65 1.32 1.65 1.32 1.285 1.38 1.285 1.38 1.65 2.035 1.65 2.035 1.25 2.095 1.25 2.095 1.65 2.435 1.65 2.435 1.51 2.495 1.51 2.495 1.65 3.49 1.65 3.49 1.54 3.61 1.54 3.61 1.65 3.96 1.65 3.96 1.38 4.08 1.38 4.08 1.44 4.02 1.44 4.02 1.65 5.135 1.65 5.135 1.51 5.195 1.51 5.195 1.65 5.88 1.65 5.88 1.51 5.94 1.51 5.94 1.65 6.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 0.06 6.04 0.06 6.04 0.17 5.92 0.17 5.92 0.06 5.135 0.06 5.135 0.5 5.075 0.5 5.075 0.06 3.68 0.06 3.68 0.17 3.56 0.17 3.56 0.06 2.55 0.06 2.55 0.26 2.43 0.26 2.43 0.2 2.49 0.2 2.49 0.06 1.35 0.06 1.35 0.47 1.29 0.47 1.29 0.06 0.915 0.06 0.915 0.47 0.855 0.47 0.855 0.06 0.505 0.06 0.505 0.47 0.445 0.47 0.445 0.06 0 0.06 0 -0.06 6.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.3 0.89 6.195 0.89 6.195 1.04 6.135 1.04 6.135 0.83 6.24 0.83 6.24 0.5 6.185 0.5 6.185 0.335 5.375 0.335 5.375 0.825 5.315 0.825 5.315 0.275 5.62 0.275 5.62 0.16 5.74 0.16 5.74 0.275 6.245 0.275 6.245 0.44 6.3 0.44 ;
      POLYGON 5.7 0.495 5.535 0.495 5.535 1.185 4.68 1.185 4.68 1.035 4.6 1.035 4.6 0.9 4.54 0.9 4.54 0.64 4.38 0.64 4.38 0.52 4.44 0.52 4.44 0.58 4.6 0.58 4.6 0.84 4.66 0.84 4.66 0.975 4.74 0.975 4.74 1.125 5.475 1.125 5.475 0.435 5.7 0.435 ;
      POLYGON 5.035 1.345 4.425 1.345 4.425 1.28 4.325 1.28 4.325 1.34 4.265 1.34 4.265 1.28 3.1 1.28 3.1 0.79 3.03 0.79 3.03 0.275 2.71 0.275 2.71 0.42 1.8 0.42 1.8 0.99 1.68 0.99 1.68 0.93 1.74 0.93 1.74 0.36 2.65 0.36 2.65 0.215 3.09 0.215 3.09 0.73 3.16 0.73 3.16 1.22 4.485 1.22 4.485 1.285 5.035 1.285 ;
      POLYGON 4.96 1.01 4.84 1.01 4.84 0.95 4.87 0.95 4.87 0.68 4.76 0.68 4.76 0.74 4.7 0.74 4.7 0.405 3.19 0.405 3.19 0.345 4.76 0.345 4.76 0.62 4.87 0.62 4.87 0.405 4.93 0.405 4.93 0.95 4.96 0.95 ;
      POLYGON 4.455 1.12 4.395 1.12 4.395 1.06 4.38 1.06 4.38 0.94 3.54 0.94 3.54 0.9 3.48 0.9 3.48 0.84 3.6 0.84 3.6 0.88 4.16 0.88 4.16 0.52 4.22 0.52 4.22 0.88 4.44 0.88 4.44 1 4.455 1 ;
      RECT 3.725 1.04 4.28 1.12 ;
      POLYGON 3.945 0.78 3.825 0.78 3.825 0.74 3.38 0.74 3.38 1.06 3.26 1.06 3.26 1 3.32 1 3.32 0.61 3.26 0.61 3.26 0.55 3.38 0.55 3.38 0.68 3.885 0.68 3.885 0.72 3.945 0.72 ;
      POLYGON 3 1.09 2.94 1.09 2.94 0.95 2.81 0.95 2.81 0.74 2.285 0.74 2.285 0.8 2.165 0.8 2.165 0.74 2.225 0.74 2.225 0.68 2.81 0.68 2.81 0.55 2.93 0.55 2.93 0.61 2.87 0.61 2.87 0.89 3 0.89 ;
      POLYGON 2.68 1.355 2.62 1.355 2.62 1.28 2.27 1.28 2.27 1.055 2.065 1.055 2.065 1.15 0.255 1.15 0.255 0.73 0.315 0.73 0.315 1.09 0.895 1.09 0.895 0.74 0.955 0.74 0.955 1.09 1.275 1.09 1.275 0.73 1.335 0.73 1.335 1.09 2.005 1.09 2.005 0.58 2.065 0.58 2.065 0.52 2.125 0.52 2.125 0.64 2.065 0.64 2.065 0.995 2.33 0.995 2.33 1.22 2.68 1.22 ;
      POLYGON 0.55 0.78 0.49 0.78 0.49 0.63 0.155 0.63 0.155 1.02 0.095 1.02 0.095 0.49 0.24 0.49 0.24 0.57 0.55 0.57 ;
  END
END SDFFRX2

MACRO SDFFRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRX4 0 0 ;
  SIZE 7.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2029 LAYER Metal1 ;
    ANTENNADIFFAREA 4.8956 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4554 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.2290295 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 71.0869565 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.19 0.545 6.72 0.545 6.72 0.79 6.74 0.79 6.74 0.95 7.17 0.95 7.17 1.34 7.11 1.34 7.11 1.01 6.76 1.01 6.76 1.34 6.66 1.34 6.66 0.545 6.6 0.545 6.6 0.485 7.19 0.485 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.2029 LAYER Metal1 ;
    ANTENNADIFFAREA 4.8956 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4554 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.2290295 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 71.0869565 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.35 1.34 6.29 1.34 6.29 1.01 5.94 1.01 5.94 1.34 5.86 1.34 5.86 0.545 5.66 0.545 5.66 0.485 6.25 0.485 6.25 0.545 5.92 0.545 5.92 0.79 5.94 0.79 5.94 0.95 6.35 0.95 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06255 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 15.7793765 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.41 0.76 5.35 0.76 5.35 0.705 4.665 0.705 4.665 0.645 4.725 0.645 4.725 0.45 4.41 0.45 4.41 0.355 3.765 0.355 3.765 0.865 3.225 0.865 3.225 0.805 3.705 0.805 3.705 0.705 3.635 0.705 3.635 0.625 3.705 0.625 3.705 0.295 4.47 0.295 4.47 0.39 4.785 0.39 4.785 0.64 5.41 0.64 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.46 0.6 1.54 1.1 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.6 1.34 1.1 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.68 1.1 0.46 1.1 0.46 0.74 0.54 0.74 0.54 0.79 0.68 0.79 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 21.85185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.16 1.1 1.1 1.1 1.1 0.315 0.6 0.315 0.6 0.58 0.695 0.58 0.695 0.625 0.755 0.625 0.755 0.685 0.635 0.685 0.635 0.64 0.34 0.64 0.34 0.73 0.26 0.73 0.26 0.6 0.28 0.6 0.28 0.58 0.54 0.58 0.54 0.255 1.16 0.255 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.8 1.77 0 1.77 0 1.65 0.475 1.65 0.475 1.36 0.535 1.36 0.535 1.65 1.335 1.65 1.335 1.36 1.395 1.36 1.395 1.65 1.975 1.65 1.975 1.285 2.035 1.285 2.035 1.65 2.79 1.65 2.79 1.54 2.91 1.54 2.91 1.65 3.57 1.65 3.57 1.55 3.51 1.55 3.51 1.49 3.63 1.49 3.63 1.65 4.41 1.65 4.41 1.125 4.47 1.125 4.47 1.65 4.94 1.65 4.94 1.22 5 1.22 5 1.65 5.675 1.65 5.675 0.95 5.735 0.95 5.735 1.65 6.085 1.65 6.085 1.11 6.145 1.11 6.145 1.65 6.495 1.65 6.495 0.95 6.555 0.95 6.555 1.65 6.905 1.65 6.905 1.11 6.965 1.11 6.965 1.65 7.345 1.65 7.345 1.02 7.405 1.02 7.405 1.65 7.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.8 0.06 7.425 0.06 7.425 0.17 7.305 0.17 7.305 0.06 6.955 0.06 6.955 0.17 6.835 0.17 6.835 0.06 6.485 0.06 6.485 0.17 6.365 0.17 6.365 0.06 6.015 0.06 6.015 0.17 5.895 0.17 5.895 0.06 5.545 0.06 5.545 0.17 5.425 0.17 5.425 0.06 4.63 0.06 4.63 0.16 4.69 0.16 4.69 0.22 4.57 0.22 4.57 0.06 3.605 0.06 3.605 0.52 3.485 0.52 3.485 0.46 3.545 0.46 3.545 0.06 1.885 0.06 1.885 0.635 1.825 0.635 1.825 0.06 1.36 0.06 1.36 0.48 1.3 0.48 1.3 0.06 0.415 0.06 0.415 0.48 0.355 0.48 0.355 0.06 0 0.06 0 -0.06 7.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.65 1.34 7.56 1.34 7.56 0.92 7.27 0.92 7.27 0.78 7.33 0.78 7.33 0.86 7.59 0.86 7.59 0.455 7.65 0.455 ;
      POLYGON 7.49 0.76 7.43 0.76 7.43 0.385 6.41 0.385 6.41 0.665 6.39 0.665 6.39 0.735 6.33 0.735 6.33 0.615 6.35 0.615 6.35 0.385 5.135 0.385 5.135 0.49 5.075 0.49 5.075 0.325 7.49 0.325 ;
      POLYGON 5.575 1.025 5.34 1.025 5.34 1.34 5.28 1.34 5.28 1.025 4.795 1.025 4.795 1.34 4.735 1.34 4.735 1.025 4.345 1.025 4.345 0.87 4.405 0.87 4.405 0.965 5.515 0.965 5.515 0.78 5.575 0.78 ;
      POLYGON 4.955 0.865 4.505 0.865 4.505 0.61 4.085 0.61 4.085 1.185 3.965 1.185 3.965 1.125 4.025 1.125 4.025 0.55 4.07 0.55 4.07 0.455 4.13 0.455 4.13 0.55 4.565 0.55 4.565 0.805 4.955 0.805 ;
      POLYGON 4.305 0.77 4.245 0.77 4.245 1.375 3.41 1.375 3.41 1.405 3.01 1.405 3.01 1.365 2.66 1.365 2.66 1.31 2.135 1.31 2.135 1.25 2.66 1.25 2.66 1.165 2.72 1.165 2.72 1.305 3.07 1.305 3.07 1.345 3.35 1.345 3.35 1.315 4.185 1.315 4.185 0.71 4.305 0.71 ;
      POLYGON 3.925 1.025 3.865 1.025 3.865 1.12 3.745 1.12 3.745 1.025 3.065 1.025 3.065 0.87 3.125 0.87 3.125 0.965 3.865 0.965 3.865 0.455 3.925 0.455 ;
      POLYGON 3.535 0.705 2.85 0.705 2.85 0.895 2.725 0.895 2.725 1.005 2.645 1.005 2.645 1.065 2.585 1.065 2.585 0.945 2.665 0.945 2.665 0.835 2.79 0.835 2.79 0.455 2.85 0.455 2.85 0.645 3.535 0.645 ;
      POLYGON 3.445 0.285 2.345 0.285 2.345 0.625 2.405 0.625 2.405 0.685 2.285 0.685 2.285 0.63 2.185 0.63 2.185 0.99 2.065 0.99 2.065 0.93 2.125 0.93 2.125 0.63 2.065 0.63 2.065 0.57 2.285 0.57 2.285 0.225 3.445 0.225 ;
      POLYGON 3.25 1.245 3.17 1.245 3.17 1.205 2.825 1.205 2.825 0.995 2.905 0.995 2.905 1.125 3.25 1.125 ;
      POLYGON 2.645 0.685 2.565 0.685 2.565 0.845 2.44 0.845 2.44 1.15 1.875 1.15 1.875 1.545 1.495 1.545 1.495 1.26 1 1.26 1 1.385 0.94 1.385 0.94 0.475 0.7 0.475 0.7 0.415 1 0.415 1 1.2 1.555 1.2 1.555 1.485 1.815 1.485 1.815 1.09 2.38 1.09 2.38 0.785 2.505 0.785 2.505 0.625 2.585 0.625 2.585 0.455 2.645 0.455 ;
      POLYGON 2.025 0.795 1.715 0.795 1.715 1.385 1.655 1.385 1.655 0.5 1.54 0.5 1.54 0.38 1.6 0.38 1.6 0.44 1.715 0.44 1.715 0.735 2.025 0.735 ;
      POLYGON 0.84 1.26 0.33 1.26 0.33 1.385 0.27 1.385 0.27 1.26 0.1 1.26 0.1 0.455 0.12 0.455 0.12 0.385 0.18 0.385 0.18 0.505 0.16 0.505 0.16 1.2 0.78 1.2 0.78 1.105 0.84 1.105 ;
  END
END SDFFRX4

MACRO SDFFRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFRXL 0 0 ;
  SIZE 6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.15595 LAYER Metal1 ;
    ANTENNADIFFAREA 3.28615 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2106 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.9855175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 114.84330475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 1.385 0.86 1.385 0.86 0.47 0.92 0.47 0.92 0.98 0.94 0.98 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.15595 LAYER Metal1 ;
    ANTENNADIFFAREA 3.28615 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2106 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.9855175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 114.84330475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.285 1.02 0.205 1.02 0.205 0.73 0.06 0.73 0.06 0.6 0.205 0.6 0.205 0.54 0.285 0.54 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 16.52777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.765 0.705 5.635 0.705 5.635 0.525 5.13 0.525 5.13 0.725 5.07 0.725 5.07 0.525 4.865 0.525 4.865 0.91 4.805 0.91 4.805 0.465 5.695 0.465 5.695 0.625 5.765 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.535 0.9 5.23 0.9 5.23 0.625 5.365 0.625 5.365 0.82 5.535 0.82 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.545 0.87 4.54 0.87 4.54 0.99 4.46 0.99 4.46 0.79 4.465 0.79 4.465 0.495 4.545 0.495 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.084 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 2.5925925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 32.4074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.11 0.9 1.765 0.9 1.765 0.92 1.635 0.92 1.635 0.815 1.765 0.815 1.765 0.82 2.11 0.82 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.21 1.085 1.14 1.085 1.14 1.26 1.06 1.26 1.06 0.98 1.13 0.98 1.13 0.83 1.21 0.83 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 1.77 0 1.77 0 1.65 0.46 1.65 0.46 0.995 0.52 0.995 0.52 1.65 1.085 1.65 1.085 1.36 1.145 1.36 1.145 1.65 1.55 1.65 1.55 1.35 1.61 1.35 1.61 1.65 1.99 1.65 1.99 1.54 2.11 1.54 2.11 1.65 2.95 1.65 2.95 1.54 3.07 1.54 3.07 1.65 3.38 1.65 3.38 1.51 3.44 1.51 3.44 1.65 4.495 1.65 4.495 1.51 4.555 1.51 4.555 1.65 5.325 1.65 5.325 1.16 5.385 1.16 5.385 1.65 6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 0.06 5.355 0.06 5.355 0.305 5.415 0.305 5.415 0.365 5.295 0.365 5.295 0.06 4.515 0.06 4.515 0.395 4.455 0.395 4.455 0.06 3.17 0.06 3.17 0.17 3.05 0.17 3.05 0.06 1.965 0.06 1.965 0.335 2.025 0.335 2.025 0.395 1.905 0.395 1.905 0.06 1.05 0.06 1.05 0.2 0.99 0.2 0.99 0.06 0.52 0.06 0.52 0.2 0.46 0.2 0.46 0.06 0 0.06 0 -0.06 6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.925 1.06 5.77 1.06 5.77 1.185 5.71 1.185 5.71 1.06 5.065 1.06 5.065 0.995 4.985 0.995 4.985 0.935 5.125 0.935 5.125 1 5.865 1 5.865 0.365 5.68 0.365 5.68 0.305 5.925 0.305 ;
      POLYGON 5.085 0.365 4.705 0.365 4.705 1.095 4.965 1.095 4.965 1.155 4.705 1.155 4.705 1.315 3.995 1.315 3.995 0.845 3.9 0.845 3.9 0.46 3.96 0.46 3.96 0.785 4.055 0.785 4.055 1.255 4.645 1.255 4.645 0.305 5.085 0.305 ;
      POLYGON 4.395 1.475 3.715 1.475 3.715 1.285 3.33 1.285 3.33 1.25 1.37 1.25 1.37 1.385 1.31 1.385 1.31 0.47 1.37 0.47 1.37 1.19 2.21 1.19 2.21 0.66 2.27 0.66 2.27 1.19 2.59 1.19 2.59 0.88 2.53 0.88 2.53 0.82 2.65 0.82 2.65 1.19 3.39 1.19 3.39 1.225 3.715 1.225 3.715 1.165 3.775 1.165 3.775 1.415 4.395 1.415 ;
      POLYGON 4.35 1.155 4.23 1.155 4.23 0.42 4.13 0.42 4.13 0.685 4.07 0.685 4.07 0.335 3.5 0.335 3.5 0.39 2.715 0.39 2.715 0.65 2.81 0.65 2.81 0.77 2.75 0.77 2.75 0.71 2.655 0.71 2.655 0.33 3.44 0.33 3.44 0.275 4.13 0.275 4.13 0.36 4.23 0.36 4.23 0.3 4.29 0.3 4.29 1.095 4.35 1.095 ;
      POLYGON 3.85 1.065 3.79 1.065 3.79 1.005 3.74 1.005 3.74 0.87 3.07 0.87 3.07 0.66 3.13 0.66 3.13 0.81 3.6 0.81 3.6 0.46 3.66 0.46 3.66 0.81 3.8 0.81 3.8 0.945 3.85 0.945 ;
      POLYGON 3.64 1.09 3.18 1.09 3.18 1.01 3.56 1.01 3.56 0.97 3.64 0.97 ;
      POLYGON 3.445 0.71 3.23 0.71 3.23 0.55 2.97 0.55 2.97 1.04 2.785 1.04 2.785 0.98 2.91 0.98 2.91 0.55 2.815 0.55 2.815 0.49 3.29 0.49 3.29 0.65 3.445 0.65 ;
      RECT 1.83 1.35 3.23 1.41 ;
      POLYGON 2.49 1.04 2.37 1.04 2.37 0.555 1.69 0.555 1.69 0.36 1.63 0.36 1.63 0.3 1.75 0.3 1.75 0.495 2.37 0.495 2.37 0.435 2.43 0.435 2.43 0.98 2.49 0.98 ;
      POLYGON 2.11 0.72 1.865 0.72 1.865 0.715 1.535 0.715 1.535 1.02 1.875 1.02 1.875 1.08 1.475 1.08 1.475 0.52 1.47 0.52 1.47 0.37 1.21 0.37 1.21 0.73 1.02 0.73 1.02 0.67 1.15 0.67 1.15 0.31 1.53 0.31 1.53 0.46 1.57 0.46 1.57 0.655 1.9 0.655 1.9 0.66 2.11 0.66 ;
      POLYGON 0.755 1.02 0.675 1.02 0.675 0.79 0.385 0.79 0.385 0.71 0.66 0.71 0.66 0.54 0.74 0.54 0.74 0.71 0.755 0.71 ;
  END
END SDFFRXL

MACRO SDFFSHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSHQX1 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.44285 LAYER Metal1 ;
    ANTENNADIFFAREA 3.80145 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2601 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.23663975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 102.4913495 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 0.92 0.66 0.92 0.66 0.87 0.56 0.87 0.56 1.02 0.48 1.02 0.48 0.57 0.6 0.57 0.6 0.65 0.56 0.65 0.56 0.79 0.74 0.79 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.8646865 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.16 0.73 6.06 0.73 6.06 0.715 5.25 0.715 5.25 0.635 6.06 0.635 6.06 0.6 6.14 0.6 6.14 0.61 6.16 0.61 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.905 1.025 5.825 1.025 5.825 0.935 5.535 0.935 5.535 0.815 5.905 0.815 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.30769225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.56 0.625 4.83 0.775 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.83 0.955 4.66 0.955 4.66 1.01 4.385 1.01 4.385 0.875 4.83 0.875 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.14239475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.505 0.975 2.445 0.975 2.445 1.18 2.05 1.18 2.05 1.28 1.565 1.28 1.565 1.295 1.08 1.295 1.08 1.11 1.06 1.11 1.06 0.98 1.08 0.98 1.08 0.875 1.14 0.875 1.14 1.235 1.505 1.235 1.505 1.22 1.99 1.22 1.99 1.12 2.385 1.12 2.385 0.915 2.505 0.915 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 1.77 0 1.77 0 1.65 0.24 1.65 0.24 0.92 0.3 0.92 0.3 1.65 1.05 1.65 1.05 1.54 1.17 1.54 1.17 1.65 1.52 1.65 1.52 1.54 1.64 1.54 1.64 1.65 2.31 1.65 2.31 1.54 2.43 1.54 2.43 1.65 2.815 1.65 2.815 1.54 2.935 1.54 2.935 1.65 4.065 1.65 4.065 0.995 4.125 0.995 4.125 1.65 4.74 1.65 4.74 1.11 4.8 1.11 4.8 1.65 5.62 1.65 5.62 1.285 5.68 1.285 5.68 1.65 6.27 1.65 6.27 1.175 6.33 1.175 6.33 1.65 6.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 0.06 6.3 0.06 6.3 0.53 6.24 0.53 6.24 0.06 5.585 0.06 5.585 0.375 5.525 0.375 5.525 0.06 4.83 0.06 4.83 0.345 4.71 0.345 4.71 0.285 4.77 0.285 4.77 0.06 4.055 0.06 4.055 0.17 3.935 0.17 3.935 0.06 3.04 0.06 3.04 0.48 2.98 0.48 2.98 0.06 2.38 0.06 2.38 0.28 2.32 0.28 2.32 0.06 1.14 0.06 1.14 0.395 1.2 0.395 1.2 0.455 1.08 0.455 1.08 0.06 0.16 0.06 0.16 0.43 0.22 0.43 0.22 0.49 0.1 0.49 0.1 0.06 0 0.06 0 -0.06 6.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.125 1.085 6.065 1.085 6.065 1.185 5.375 1.185 5.375 0.875 5.09 0.875 5.09 0.475 5.685 0.475 5.685 0.44 6.06 0.44 6.06 0.5 5.745 0.5 5.745 0.535 5.15 0.535 5.15 0.815 5.435 0.815 5.435 1.125 6.005 1.125 6.005 1.025 6.125 1.025 ;
      POLYGON 5.37 1.405 5.31 1.405 5.31 1.345 5.215 1.345 5.215 1.035 4.93 1.035 4.93 0.505 4.55 0.505 4.55 0.325 4.17 0.325 4.17 0.33 3.68 0.33 3.68 1.22 3.74 1.22 3.74 1.28 3.62 1.28 3.62 0.27 4.11 0.27 4.11 0.265 4.61 0.265 4.61 0.445 4.93 0.445 4.93 0.315 5.245 0.315 5.245 0.375 4.99 0.375 4.99 0.975 5.275 0.975 5.275 1.285 5.37 1.285 ;
      POLYGON 4.565 1.23 4.505 1.23 4.505 1.17 4.225 1.17 4.225 0.75 3.97 0.75 3.97 0.69 4.225 0.69 4.225 0.425 4.45 0.425 4.45 0.485 4.285 0.485 4.285 1.11 4.565 1.11 ;
      POLYGON 3.91 0.585 3.85 0.585 3.85 0.9 3.9 0.9 3.9 1.44 1.85 1.44 1.85 1.38 3.46 1.38 3.46 0.91 3.52 0.91 3.52 1.38 3.84 1.38 3.84 0.96 3.79 0.96 3.79 0.525 3.91 0.525 ;
      POLYGON 3.52 0.725 3.46 0.725 3.46 0.345 3.2 0.345 3.2 0.97 3.14 0.97 3.14 0.64 2.82 0.64 2.82 0.44 2.22 0.44 2.22 0.64 2.16 0.64 2.16 0.36 1.62 0.36 1.62 0.62 1.63 0.62 1.63 0.74 1.56 0.74 1.56 0.3 2.22 0.3 2.22 0.38 2.88 0.38 2.88 0.58 3.14 0.58 3.14 0.285 3.52 0.285 ;
      POLYGON 3.36 1.19 3.3 1.19 3.3 1.13 2.765 1.13 2.765 0.9 2.825 0.9 2.825 1.07 3.3 1.07 3.3 0.445 3.36 0.445 ;
      POLYGON 3.04 0.8 2.665 0.8 2.665 1.16 2.545 1.16 2.545 1.1 2.605 1.1 2.605 0.8 2.22 0.8 2.22 1.02 2.16 1.02 2.16 0.8 2 0.8 2 0.54 1.94 0.54 1.94 0.48 2.06 0.48 2.06 0.74 2.66 0.74 2.66 0.54 2.72 0.54 2.72 0.74 3.04 0.74 ;
      POLYGON 2.015 1.02 1.955 1.02 1.955 0.96 1.84 0.96 1.84 0.9 1.24 0.9 1.24 0.775 1.015 0.775 1.015 0.715 1.3 0.715 1.3 0.84 1.78 0.84 1.78 0.52 1.72 0.52 1.72 0.46 1.84 0.46 1.84 0.84 1.9 0.84 1.9 0.9 2.015 0.9 ;
      POLYGON 1.74 1.12 1.405 1.12 1.405 1.135 1.285 1.135 1.285 1.055 1.325 1.055 1.325 1.04 1.66 1.04 1.66 1 1.74 1 ;
      POLYGON 1.46 0.73 1.4 0.73 1.4 0.615 0.915 0.615 0.915 1.08 0.905 1.08 0.905 1.165 0.845 1.165 0.845 1.02 0.855 1.02 0.855 0.47 0.38 0.47 0.38 0.82 0.32 0.82 0.32 0.41 0.965 0.41 0.965 0.555 1.46 0.555 ;
  END
END SDFFSHQX1

MACRO SDFFSHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSHQX2 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5541 LAYER Metal1 ;
    ANTENNADIFFAREA 3.809675 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.28935 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.28304825 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 95.81130125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.5 1.29 0.42 1.29 0.42 0.705 0.235 0.705 0.235 0.625 0.42 0.625 0.42 0.51 0.5 0.51 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.23762375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.34 0.73 6.26 0.73 6.26 0.715 5.525 0.715 5.525 0.635 6.26 0.635 6.26 0.6 6.34 0.6 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.16 0.895 5.825 0.895 5.825 0.98 5.745 0.98 5.745 0.815 6.16 0.815 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.98 0.79 4.86 0.79 4.86 0.705 4.565 0.705 4.565 0.625 4.98 0.625 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.945 0.97 4.765 0.97 4.765 1.085 4.56 1.085 4.56 0.89 4.945 0.89 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.368932 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.605 1.025 2.545 1.025 2.545 1.245 1.105 1.245 1.105 0.895 1.035 0.895 1.035 0.815 1.165 0.815 1.165 1.185 2.485 1.185 2.485 0.965 2.605 0.965 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 1.77 0 1.77 0 1.65 0.235 1.65 0.235 0.9 0.295 0.9 0.295 1.65 0.645 1.65 0.645 0.9 0.705 0.9 0.705 1.65 1.095 1.65 1.095 1.54 1.215 1.54 1.215 1.65 1.565 1.65 1.565 1.54 1.685 1.54 1.685 1.65 2.47 1.65 2.47 1.54 2.59 1.54 2.59 1.65 2.94 1.65 2.94 1.54 3.06 1.54 3.06 1.65 4.18 1.65 4.18 0.995 4.24 0.995 4.24 1.65 5.045 1.65 5.045 0.985 5.105 0.985 5.105 1.65 5.8 1.65 5.8 1.255 5.86 1.255 5.86 1.65 6.27 1.65 6.27 0.995 6.33 0.995 6.33 1.65 6.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 0.06 6.33 0.06 6.33 0.5 6.27 0.5 6.27 0.06 5.86 0.06 5.86 0.375 5.8 0.375 5.8 0.06 5.105 0.06 5.105 0.345 4.985 0.345 4.985 0.285 5.045 0.285 5.045 0.06 4.34 0.06 4.34 0.17 4.22 0.17 4.22 0.06 3.175 0.06 3.175 0.505 3.115 0.505 3.115 0.06 2.475 0.06 2.475 0.49 2.415 0.49 2.415 0.06 1.155 0.06 1.155 0.335 1.215 0.335 1.215 0.395 1.095 0.395 1.095 0.06 0.73 0.06 0.73 0.49 0.67 0.49 0.67 0.06 0.295 0.06 0.295 0.49 0.235 0.49 0.235 0.06 0 0.06 0 -0.06 6.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.155 1.085 6.095 1.085 6.095 1.14 5.585 1.14 5.585 0.915 5.365 0.915 5.365 0.685 5.24 0.685 5.24 0.625 5.365 0.625 5.365 0.475 5.96 0.475 5.96 0.435 6.09 0.435 6.09 0.495 6.02 0.495 6.02 0.535 5.425 0.535 5.425 0.855 5.645 0.855 5.645 1.08 6.035 1.08 6.035 1.025 6.155 1.025 ;
      POLYGON 5.485 1.375 5.425 1.375 5.425 1.075 5.205 1.075 5.205 0.845 5.08 0.845 5.08 0.505 4.825 0.505 4.825 0.325 4.505 0.325 4.505 0.33 3.875 0.33 3.875 1.215 3.755 1.215 3.755 1.095 3.815 1.095 3.815 0.27 4.445 0.27 4.445 0.265 4.885 0.265 4.885 0.445 5.205 0.445 5.205 0.315 5.425 0.315 5.425 0.375 5.265 0.375 5.265 0.505 5.14 0.505 5.14 0.785 5.265 0.785 5.265 1.015 5.485 1.015 ;
      POLYGON 4.725 0.49 4.46 0.49 4.46 1.185 4.705 1.185 4.705 1.305 4.645 1.305 4.645 1.245 4.4 1.245 4.4 0.77 4.135 0.77 4.135 0.71 4.4 0.71 4.4 0.43 4.605 0.43 4.605 0.425 4.725 0.425 ;
      POLYGON 4.105 0.61 4.035 0.61 4.035 1.375 2.705 1.375 2.705 1.405 1.845 1.405 1.845 1.345 2.645 1.345 2.645 1.315 3.595 1.315 3.595 0.935 3.655 0.935 3.655 1.315 3.975 1.315 3.975 0.55 4.105 0.55 ;
      POLYGON 3.715 0.75 3.655 0.75 3.655 0.4 3.335 0.4 3.335 0.885 3.215 0.885 3.215 0.825 3.275 0.825 3.275 0.665 2.955 0.665 2.955 0.385 2.635 0.385 2.635 0.65 2.375 0.65 2.375 0.705 2.255 0.705 2.255 0.305 1.645 0.305 1.645 0.625 1.655 0.625 1.655 0.745 1.585 0.745 1.585 0.245 2.315 0.245 2.315 0.59 2.575 0.59 2.575 0.325 3.015 0.325 3.015 0.605 3.275 0.605 3.275 0.34 3.715 0.34 ;
      POLYGON 3.555 0.56 3.495 0.56 3.495 1.215 3.435 1.215 3.435 1.045 2.865 1.045 2.865 0.925 2.925 0.925 2.925 0.985 3.435 0.985 3.435 0.5 3.555 0.5 ;
      POLYGON 3.115 0.825 2.765 0.825 2.765 1.145 2.825 1.145 2.825 1.205 2.705 1.205 2.705 0.825 2.525 0.825 2.525 0.865 2.215 0.865 2.215 1.02 2.155 1.02 2.155 0.865 2.095 0.865 2.095 0.575 1.95 0.575 1.95 0.455 2.01 0.455 2.01 0.515 2.155 0.515 2.155 0.805 2.465 0.805 2.465 0.765 2.735 0.765 2.735 0.485 2.855 0.485 2.855 0.545 2.795 0.545 2.795 0.765 3.115 0.765 ;
      POLYGON 2.01 1.085 1.95 1.085 1.95 1.025 1.935 1.025 1.935 0.905 1.265 0.905 1.265 0.715 1.035 0.715 1.035 0.655 1.325 0.655 1.325 0.845 1.755 0.845 1.755 0.525 1.745 0.525 1.745 0.405 1.805 0.405 1.805 0.465 1.815 0.465 1.815 0.845 1.995 0.845 1.995 0.965 2.01 0.965 ;
      RECT 1.33 1.005 1.835 1.085 ;
      POLYGON 1.485 0.735 1.425 0.735 1.425 0.555 0.935 0.555 0.935 1.21 0.875 1.21 0.875 0.76 0.6 0.76 0.6 0.7 0.875 0.7 0.875 0.435 0.935 0.435 0.935 0.495 1.485 0.495 ;
  END
END SDFFSHQX2

MACRO SDFFSHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSHQX4 0 0 ;
  SIZE 7.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.16171625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.98 0.705 6.94 0.705 6.94 0.73 6.86 0.73 6.86 0.715 6.025 0.715 6.025 0.655 6.86 0.655 6.86 0.6 6.94 0.6 6.94 0.645 6.98 0.645 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.76 0.895 6.395 0.895 6.395 0.95 6.315 0.95 6.315 0.815 6.76 0.815 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.545 0.895 5.465 0.895 5.465 0.705 5.235 0.705 5.235 0.625 5.545 0.625 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.305 0.895 5.035 0.895 5.035 0.685 5.015 0.685 5.015 0.605 5.135 0.605 5.135 0.815 5.305 0.815 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 16.24595475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.125 1.06 3.065 1.06 3.065 1.265 2 1.265 2 1.305 1.48 1.305 1.48 1.3 1.46 1.3 1.46 1.17 1.48 1.17 1.48 0.835 1.67 0.835 1.67 0.895 1.54 0.895 1.54 1.245 1.94 1.245 1.94 1.205 3.005 1.205 3.005 1 3.125 1 ;
    END
  END SN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.88455 LAYER Metal1 ;
    ANTENNADIFFAREA 4.407225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.371025 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.46977975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 81.9567415 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.905 0.66 0.86 0.66 0.86 0.91 0.905 0.91 0.905 1.355 0.845 1.355 0.845 0.97 0.8 0.97 0.8 0.705 0.54 0.705 0.54 0.73 0.495 0.73 0.495 1.355 0.435 1.355 0.435 0.54 0.495 0.54 0.495 0.6 0.54 0.6 0.54 0.645 0.8 0.645 0.8 0.6 0.845 0.6 0.845 0.54 0.905 0.54 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 1.77 0 1.77 0 1.65 0.23 1.65 0.23 0.965 0.29 0.965 0.29 1.65 0.64 1.65 0.64 0.965 0.7 0.965 0.7 1.65 1.085 1.65 1.085 1.51 1.145 1.51 1.145 1.65 1.57 1.65 1.57 1.51 1.63 1.51 1.63 1.65 2.1 1.65 2.1 1.365 2.16 1.365 2.16 1.65 2.99 1.65 2.99 1.54 3.11 1.54 3.11 1.65 3.46 1.65 3.46 1.54 3.58 1.54 3.58 1.65 4.695 1.65 4.695 0.995 4.755 0.995 4.755 1.65 5.545 1.65 5.545 0.995 5.605 0.995 5.605 1.65 6.39 1.65 6.39 1.255 6.45 1.255 6.45 1.65 6.955 1.65 6.955 0.995 7.015 0.995 7.015 1.65 7.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 0.06 7.015 0.06 7.015 0.5 6.955 0.5 6.955 0.06 6.36 0.06 6.36 0.395 6.3 0.395 6.3 0.06 5.605 0.06 5.605 0.365 5.485 0.365 5.485 0.305 5.545 0.305 5.545 0.06 4.94 0.06 4.94 0.17 4.82 0.17 4.82 0.06 3.69 0.06 3.69 0.565 3.63 0.565 3.63 0.06 2.99 0.06 2.99 0.565 2.93 0.565 2.93 0.06 1.6 0.06 1.6 0.355 1.66 0.355 1.66 0.415 1.54 0.415 1.54 0.06 1.11 0.06 1.11 0.52 1.05 0.52 1.05 0.06 0.7 0.06 0.7 0.52 0.64 0.52 0.64 0.06 0.29 0.06 0.29 0.52 0.23 0.52 0.23 0.06 0 0.06 0 -0.06 7.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.84 1.085 6.78 1.085 6.78 1.11 5.865 1.11 5.865 0.685 5.805 0.685 5.805 0.625 5.865 0.625 5.865 0.495 6.655 0.495 6.655 0.435 6.775 0.435 6.775 0.495 6.715 0.495 6.715 0.555 5.925 0.555 5.925 0.855 6.215 0.855 6.215 0.915 5.925 0.915 5.925 1.05 6.72 1.05 6.72 1.025 6.84 1.025 ;
      POLYGON 6.14 1.33 6.08 1.33 6.08 1.27 5.705 1.27 5.705 0.895 5.645 0.895 5.645 0.525 5.325 0.525 5.325 0.345 4.39 0.345 4.39 1.215 4.33 1.215 4.33 1.275 4.27 1.275 4.27 1.155 4.33 1.155 4.33 0.285 5.385 0.285 5.385 0.465 5.705 0.465 5.705 0.335 5.99 0.335 5.99 0.395 5.765 0.395 5.765 0.525 5.705 0.525 5.705 0.835 5.765 0.835 5.765 1.21 6.14 1.21 ;
      POLYGON 5.3 1.115 5.24 1.115 5.24 1.055 4.855 1.055 4.855 0.79 4.65 0.79 4.65 0.73 4.855 0.73 4.855 0.445 5.225 0.445 5.225 0.505 4.915 0.505 4.915 0.995 5.3 0.995 ;
      POLYGON 4.705 0.63 4.55 0.63 4.55 1.435 3.79 1.435 3.79 1.425 2.38 1.425 2.38 1.365 3.85 1.365 3.85 1.375 4.11 1.375 4.11 0.995 4.17 0.995 4.17 1.375 4.49 1.375 4.49 0.57 4.705 0.57 ;
      POLYGON 4.23 0.81 4.17 0.81 4.17 0.46 3.85 0.46 3.85 0.945 3.73 0.945 3.73 0.885 3.79 0.885 3.79 0.725 3.47 0.725 3.47 0.46 3.15 0.46 3.15 0.725 2.74 0.725 2.74 0.415 2.15 0.415 2.15 0.685 2.21 0.685 2.21 0.745 2.09 0.745 2.09 0.355 2.8 0.355 2.8 0.665 3.09 0.665 3.09 0.4 3.53 0.4 3.53 0.665 3.79 0.665 3.79 0.4 4.23 0.4 ;
      POLYGON 4.07 0.62 4.01 0.62 4.01 1.275 3.95 1.275 3.95 1.105 3.385 1.105 3.385 0.985 3.445 0.985 3.445 1.045 3.95 1.045 3.95 0.56 4.07 0.56 ;
      POLYGON 3.63 0.885 3.285 0.885 3.285 1.205 3.345 1.205 3.345 1.265 3.225 1.265 3.225 0.885 2.75 0.885 2.75 1.02 2.69 1.02 2.69 0.885 2.58 0.885 2.58 0.575 2.47 0.575 2.47 0.515 2.64 0.515 2.64 0.825 3.31 0.825 3.31 0.62 3.25 0.62 3.25 0.56 3.37 0.56 3.37 0.825 3.63 0.825 ;
      POLYGON 2.545 1.105 2.485 1.105 2.485 1.045 2.42 1.045 2.42 0.925 1.77 0.925 1.77 0.735 1.37 0.735 1.37 0.675 1.83 0.675 1.83 0.865 2.31 0.865 2.31 0.575 2.25 0.575 2.25 0.515 2.37 0.515 2.37 0.865 2.48 0.865 2.48 0.985 2.545 0.985 ;
      POLYGON 2.32 1.105 1.84 1.105 1.84 1.145 1.76 1.145 1.76 1.025 2.32 1.025 ;
      POLYGON 1.99 0.765 1.93 0.765 1.93 0.575 1.27 0.575 1.27 0.965 1.36 0.965 1.36 1.275 1.3 1.275 1.3 1.025 1.21 1.025 1.21 0.815 0.96 0.815 0.96 0.755 1.21 0.755 1.21 0.515 1.3 0.515 1.3 0.455 1.36 0.455 1.36 0.515 1.99 0.515 ;
  END
END SDFFSHQX4

MACRO SDFFSHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSHQX8 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.4542 LAYER Metal1 ;
    ANTENNADIFFAREA 5.21655 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.528525 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.42760525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 66.17851575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.68 0.99 1.565 0.99 1.565 1.05 1.505 1.05 1.505 0.99 1.155 0.99 1.155 1.345 1.095 1.345 1.095 0.73 1.06 0.73 1.06 0.66 0.745 0.66 0.745 1.345 0.685 1.345 0.685 0.66 0.335 0.66 0.335 1.345 0.275 1.345 0.275 0.54 0.335 0.54 0.335 0.6 0.685 0.6 0.685 0.54 0.745 0.54 0.745 0.6 1.095 0.6 1.095 0.54 1.155 0.54 1.155 0.93 1.62 0.93 1.62 0.54 1.68 0.54 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.16171625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.94 0.92 7.86 0.92 7.86 0.79 7.045 0.79 7.045 0.73 7.92 0.73 7.92 0.79 7.94 0.79 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.32 0.945 7.76 1.085 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.61 0.89 6.365 0.89 6.365 0.905 6.235 0.905 6.235 0.7 6.365 0.7 6.365 0.81 6.61 0.81 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.265 1.085 6.035 1.085 6.035 0.835 6.015 0.835 6.015 0.755 6.135 0.755 6.135 1.005 6.265 1.005 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.724919 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.94 1.01 3.835 1.01 3.835 1.28 3.575 1.28 3.575 1.35 2.505 1.35 2.505 1.085 2.435 1.085 2.435 1.005 2.505 1.005 2.505 0.93 2.575 0.93 2.575 1.05 2.565 1.05 2.565 1.29 3.515 1.29 3.515 1.22 3.775 1.22 3.775 0.95 3.94 0.95 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.9 0.13 0.9 0.13 1.65 0.48 1.65 0.48 0.9 0.54 0.9 0.54 1.65 0.89 1.65 0.89 0.9 0.95 0.9 0.95 1.65 1.3 1.65 1.3 1.09 1.36 1.09 1.36 1.65 1.95 1.65 1.95 0.9 2.01 0.9 2.01 1.65 2.36 1.65 2.36 1.45 2.48 1.45 2.48 1.51 2.42 1.51 2.42 1.65 2.9 1.65 2.9 1.45 3.02 1.45 3.02 1.51 2.96 1.51 2.96 1.65 3.835 1.65 3.835 1.54 3.955 1.54 3.955 1.65 4.305 1.65 4.305 1.54 4.425 1.54 4.425 1.65 5.495 1.65 5.495 0.995 5.555 0.995 5.555 1.65 6.535 1.65 6.535 1.085 6.595 1.085 6.595 1.65 7.425 1.65 7.425 1.355 7.485 1.355 7.485 1.65 7.87 1.65 7.87 1.345 7.93 1.345 7.93 1.65 8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 0.06 7.86 0.06 7.86 0.2 7.8 0.2 7.8 0.06 7.38 0.06 7.38 0.47 7.32 0.47 7.32 0.06 6.625 0.06 6.625 0.44 6.505 0.44 6.505 0.38 6.565 0.38 6.565 0.06 5.75 0.06 5.75 0.335 5.63 0.335 5.63 0.275 5.69 0.275 5.69 0.06 4.44 0.06 4.44 0.52 4.38 0.52 4.38 0.06 3.74 0.06 3.74 0.475 3.68 0.475 3.68 0.06 2.515 0.06 2.515 0.43 2.575 0.43 2.575 0.49 2.455 0.49 2.455 0.06 2.115 0.06 2.115 0.52 2.055 0.52 2.055 0.06 1.36 0.06 1.36 0.485 1.3 0.485 1.3 0.06 0.95 0.06 0.95 0.485 0.89 0.485 0.89 0.06 0.54 0.06 0.54 0.485 0.48 0.485 0.48 0.06 0.13 0.06 0.13 0.485 0.07 0.485 0.07 0.06 0 0.06 0 -0.06 8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.725 0.63 6.945 0.63 6.945 0.89 7.22 0.89 7.22 1.185 7.725 1.185 7.725 1.245 7.16 1.245 7.16 0.95 6.87 0.95 6.87 0.78 6.885 0.78 6.885 0.57 7.725 0.57 ;
      POLYGON 7.175 1.465 7.115 1.465 7.115 1.405 7 1.405 7 1.11 6.71 1.11 6.71 0.6 6.345 0.6 6.345 0.42 5.91 0.42 5.91 0.495 5.47 0.495 5.47 0.335 5.14 0.335 5.14 1.2 5.08 1.2 5.08 0.275 5.53 0.275 5.53 0.435 5.85 0.435 5.85 0.36 6.405 0.36 6.405 0.54 6.725 0.54 6.725 0.41 7.1 0.41 7.1 0.47 6.785 0.47 6.785 0.6 6.77 0.6 6.77 1.05 7.06 1.05 7.06 1.345 7.175 1.345 ;
      POLYGON 6.13 0.655 5.915 0.655 5.915 1.185 6.1 1.185 6.1 1.305 6.04 1.305 6.04 1.245 5.855 1.245 5.855 0.655 5.4 0.655 5.4 0.595 6.01 0.595 6.01 0.52 6.13 0.52 ;
      POLYGON 5.37 0.495 5.3 0.495 5.3 0.9 5.35 0.9 5.35 1.36 3.995 1.36 3.995 1.44 3.735 1.44 3.735 1.51 3.305 1.51 3.305 1.45 3.675 1.45 3.675 1.38 3.935 1.38 3.935 1.3 4.92 1.3 4.92 0.92 4.98 0.92 4.98 1.3 5.29 1.3 5.29 0.96 5.24 0.96 5.24 0.435 5.37 0.435 ;
      POLYGON 4.98 0.765 4.92 0.765 4.92 0.36 4.6 0.36 4.6 0.62 4.66 0.62 4.66 0.98 4.6 0.98 4.6 0.68 4.22 0.68 4.22 0.37 3.9 0.37 3.9 0.635 3.64 0.635 3.64 0.69 3.52 0.69 3.52 0.41 3.055 0.41 3.055 0.73 3.065 0.73 3.065 0.85 2.995 0.85 2.995 0.35 3.58 0.35 3.58 0.575 3.84 0.575 3.84 0.31 4.28 0.31 4.28 0.62 4.54 0.62 4.54 0.3 4.98 0.3 ;
      POLYGON 4.82 1.2 4.76 1.2 4.76 1.14 4.29 1.14 4.29 1 4.2 1 4.2 0.94 4.35 0.94 4.35 1.08 4.76 1.08 4.76 0.52 4.7 0.52 4.7 0.46 4.82 0.46 ;
      POLYGON 4.5 0.84 4.1 0.84 4.1 1.11 4.19 1.11 4.19 1.17 4.04 1.17 4.04 0.85 3.675 0.85 3.675 1.02 3.615 1.02 3.615 0.85 3.36 0.85 3.36 0.54 3.42 0.54 3.42 0.79 4 0.79 4 0.47 4.12 0.47 4.12 0.53 4.06 0.53 4.06 0.78 4.5 0.78 ;
      POLYGON 3.47 1.07 3.41 1.07 3.41 1.01 2.675 1.01 2.675 0.83 2.315 0.83 2.315 0.77 2.735 0.77 2.735 0.95 3.165 0.95 3.165 0.63 3.155 0.63 3.155 0.51 3.215 0.51 3.215 0.57 3.225 0.57 3.225 0.95 3.47 0.95 ;
      RECT 2.665 1.11 3.295 1.19 ;
      POLYGON 2.895 0.82 2.835 0.82 2.835 0.67 2.215 0.67 2.215 1.29 2.155 1.29 2.155 0.68 1.85 0.68 1.85 1.135 1.805 1.135 1.805 1.195 1.745 1.195 1.745 1.075 1.79 1.075 1.79 0.44 1.52 0.44 1.52 0.83 1.46 0.83 1.46 0.38 1.85 0.38 1.85 0.4 1.91 0.4 1.91 0.62 2.175 0.62 2.175 0.61 2.26 0.61 2.26 0.54 2.32 0.54 2.32 0.61 2.895 0.61 ;
  END
END SDFFSHQX8

MACRO SDFFSRHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRHQX1 0 0 ;
  SIZE 7.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3118 LAYER Metal1 ;
    ANTENNADIFFAREA 4.627875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.30645 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.07015825 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 110.8565835 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.17 1.29 0.11 1.29 0.11 0.73 0.06 0.73 0.06 0.6 0.08 0.6 0.08 0.51 0.14 0.51 0.14 0.67 0.17 0.67 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.73267325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.565 0.705 6.885 0.705 6.885 0.905 6.825 0.905 6.825 0.645 7.39 0.645 7.39 0.625 7.565 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.61 0.895 7.34 0.895 7.34 0.98 7.205 0.98 7.205 0.81 7.235 0.81 7.235 0.805 7.34 0.805 7.34 0.815 7.61 0.815 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.12820525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.435 0.54 6.565 0.91 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.335 0.895 6.165 0.895 6.165 0.91 5.85 0.91 5.85 0.815 6.335 0.815 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 23.85113275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.28 1.385 3.58 1.385 3.58 1.22 3.26 1.22 3.26 1.355 2.4 1.355 2.4 1.005 1.48 1.005 1.48 0.92 1.46 0.92 1.46 0.79 1.54 0.79 1.54 0.945 2.46 0.945 2.46 1.295 3.2 1.295 3.2 1.16 3.64 1.16 3.64 1.325 4.28 1.325 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.92 1.26 0.92 1.26 0.91 1.025 0.91 1.025 0.655 1.105 0.655 1.105 0.79 1.34 0.79 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.8 1.77 0 1.77 0 1.65 0.315 1.65 0.315 1.06 0.375 1.06 0.375 1.65 1.16 1.65 1.16 1.24 1.1 1.24 1.1 1.18 1.22 1.18 1.22 1.65 1.96 1.65 1.96 1.265 2.08 1.265 2.08 1.325 2.02 1.325 2.02 1.65 3.42 1.65 3.42 1.38 3.36 1.38 3.36 1.32 3.48 1.32 3.48 1.65 4.38 1.65 4.38 1.295 4.5 1.295 4.5 1.355 4.44 1.355 4.44 1.65 5.85 1.65 5.85 1.17 5.91 1.17 5.91 1.65 6.575 1.65 6.575 1.24 6.635 1.24 6.635 1.65 7.27 1.65 7.27 1.24 7.33 1.24 7.33 1.65 7.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.8 0.06 7.405 0.06 7.405 0.525 7.345 0.525 7.345 0.06 6.635 0.06 6.635 0.17 6.515 0.17 6.515 0.06 5.755 0.06 5.755 0.17 5.635 0.17 5.635 0.06 4.485 0.06 4.485 0.335 4.545 0.335 4.545 0.395 4.425 0.395 4.425 0.06 1.38 0.06 1.38 0.17 1.26 0.17 1.26 0.06 0.345 0.06 0.345 0.545 0.285 0.545 0.285 0.06 0 0.06 0 -0.06 7.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.77 1.14 7.535 1.14 7.535 1.265 7.475 1.265 7.475 1.14 7.045 1.14 7.045 0.9 6.985 0.9 6.985 0.84 7.105 0.84 7.105 1.08 7.71 1.08 7.71 0.52 7.52 0.52 7.52 0.46 7.77 0.46 ;
      POLYGON 7.125 0.405 6.825 0.405 6.825 0.385 6.725 0.385 6.725 1.005 6.945 1.005 6.945 1.36 6.885 1.36 6.885 1.065 6.665 1.065 6.665 0.385 5.2 0.385 5.2 0.645 5.42 0.645 5.42 1.035 5.3 1.035 5.3 0.975 5.36 0.975 5.36 0.705 5.14 0.705 5.14 0.325 6.885 0.325 6.885 0.345 7.125 0.345 ;
      POLYGON 6.46 1.235 6.34 1.235 6.34 1.07 5.75 1.07 5.75 1.355 4.6 1.355 4.6 1.195 3.74 1.195 3.74 1.06 3.1 1.06 3.1 1.195 2.72 1.195 2.72 0.68 2.78 0.68 2.78 0.365 2.46 0.365 2.46 0.685 2.34 0.685 2.34 0.625 2.4 0.625 2.4 0.305 2.84 0.305 2.84 0.74 2.78 0.74 2.78 1.135 3.04 1.135 3.04 1 3.8 1 3.8 1.135 4.66 1.135 4.66 1.295 5.69 1.295 5.69 0.485 6.27 0.485 6.27 0.545 5.75 0.545 5.75 1.01 6.4 1.01 6.4 1.175 6.46 1.175 ;
      POLYGON 5.59 1.195 4.76 1.195 4.76 0.715 4.44 0.715 4.44 0.845 4.06 0.845 4.06 0.72 3.1 0.72 3.1 0.66 4.12 0.66 4.12 0.785 4.38 0.785 4.38 0.655 4.88 0.655 4.88 0.735 4.82 0.735 4.82 1.135 5.14 1.135 5.14 0.805 5.26 0.805 5.26 0.865 5.2 0.865 5.2 1.135 5.53 1.135 5.53 0.545 5.47 0.545 5.47 0.485 5.59 0.485 ;
      POLYGON 5.04 1.035 4.92 1.035 4.92 0.975 4.98 0.975 4.98 0.555 4.28 0.555 4.28 0.685 4.22 0.685 4.22 0.495 4.865 0.495 4.865 0.39 4.925 0.39 4.925 0.495 5.04 0.495 ;
      POLYGON 4.66 0.875 4.6 0.875 4.6 1.035 3.9 1.035 3.9 0.9 2.94 0.9 2.94 1.035 2.88 1.035 2.88 0.84 2.94 0.84 2.94 0.435 3 0.435 3 0.5 3.835 0.5 3.835 0.425 3.955 0.425 3.955 0.485 3.895 0.485 3.895 0.56 3 0.56 3 0.84 3.96 0.84 3.96 0.975 4.54 0.975 4.54 0.815 4.66 0.815 ;
      POLYGON 4.135 0.43 4.055 0.43 4.055 0.325 3.735 0.325 3.735 0.4 3.615 0.4 3.615 0.32 3.655 0.32 3.655 0.245 4.135 0.245 ;
      POLYGON 2.68 0.525 2.62 0.525 2.62 1.195 2.56 1.195 2.56 0.845 1.64 0.845 1.64 0.69 1.365 0.69 1.365 0.395 0.505 0.395 0.505 0.8 0.445 0.8 0.445 0.335 1.425 0.335 1.425 0.63 1.7 0.63 1.7 0.785 2.56 0.785 2.56 0.465 2.68 0.465 ;
      POLYGON 2.3 0.525 2.24 0.525 2.24 0.685 1.8 0.685 1.8 0.53 1.705 0.53 1.705 0.45 1.88 0.45 1.88 0.605 2.16 0.605 2.16 0.445 2.3 0.445 ;
      POLYGON 2.3 1.225 2.24 1.225 2.24 1.165 1.585 1.165 1.585 1.225 1.525 1.225 1.525 1.105 2.3 1.105 ;
      POLYGON 2.06 0.505 1.98 0.505 1.98 0.35 1.605 0.35 1.605 0.505 1.525 0.505 1.525 0.27 2.06 0.27 ;
      POLYGON 1.86 1.485 1.32 1.485 1.32 1.08 0.865 1.08 0.865 0.495 0.985 0.495 0.985 0.555 0.925 0.555 0.925 1.02 1.38 1.02 1.38 1.425 1.86 1.425 ;
      POLYGON 1.06 1.475 0.52 1.475 0.52 1.17 0.605 1.17 0.605 0.96 0.27 0.96 0.27 0.74 0.33 0.74 0.33 0.9 0.605 0.9 0.605 0.51 0.665 0.51 0.665 1.23 0.58 1.23 0.58 1.415 1.06 1.415 ;
  END
END SDFFSRHQX1

MACRO SDFFSRHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRHQX2 0 0 ;
  SIZE 8.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5362 LAYER Metal1 ;
    ANTENNADIFFAREA 4.869175 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3357 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.51266 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 106.005362 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 1.3 0.445 1.3 0.445 1.09 0.4 1.09 0.4 0.8 0.36 0.8 0.36 0.54 0.42 0.54 0.42 0.74 0.46 0.74 0.46 1.03 0.505 1.03 0.505 1.17 0.54 1.17 ;
    END
  END Q
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.4059405 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.94 0.92 7.86 0.92 7.86 0.715 7.06 0.715 7.06 0.935 7 0.935 7 0.655 7.92 0.655 7.92 0.715 7.94 0.715 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.76 1.015 7.435 1.015 7.435 0.93 7.38 0.93 7.38 0.85 7.435 0.85 7.435 0.815 7.76 0.815 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.66 0.5 6.74 1 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.56 0.895 6.215 0.895 6.215 0.815 6.48 0.815 6.48 0.66 6.56 0.66 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 24.59546925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.64 1.34 3.88 1.34 3.88 1.215 3.56 1.215 3.56 1.35 2.7 1.35 2.7 1 1.72 1 1.72 0.895 1.635 0.895 1.635 0.815 1.78 0.815 1.78 0.94 2.76 0.94 2.76 1.29 3.5 1.29 3.5 1.155 3.94 1.155 3.94 1.28 4.64 1.28 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.535 0.83 1.34 0.83 1.34 1 1.26 1 1.26 0.83 1.205 0.83 1.205 0.75 1.535 0.75 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.2 1.77 0 1.77 0 1.65 0.24 1.65 0.24 0.9 0.3 0.9 0.3 1.65 0.65 1.65 0.65 1.035 0.71 1.035 0.71 1.65 1.4 1.65 1.4 1.32 1.34 1.32 1.34 1.26 1.46 1.26 1.46 1.65 2.19 1.65 2.19 1.26 2.31 1.26 2.31 1.32 2.25 1.32 2.25 1.65 3.72 1.65 3.72 1.375 3.66 1.375 3.66 1.315 3.78 1.315 3.78 1.65 4.74 1.65 4.74 1.22 4.86 1.22 4.86 1.28 4.8 1.28 4.8 1.65 6.21 1.65 6.21 1.155 6.27 1.155 6.27 1.65 6.66 1.65 6.66 1.1 6.72 1.1 6.72 1.65 7.435 1.65 7.435 1.275 7.495 1.275 7.495 1.65 8.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.2 0.06 7.61 0.06 7.61 0.555 7.55 0.555 7.55 0.06 6.81 0.06 6.81 0.17 6.69 0.17 6.69 0.06 6.225 0.06 6.225 0.17 6.105 0.17 6.105 0.06 4.86 0.06 4.86 0.425 4.8 0.425 4.8 0.06 1.61 0.06 1.61 0.49 1.55 0.49 1.55 0.06 0.625 0.06 0.625 0.52 0.565 0.52 0.565 0.06 0.215 0.06 0.215 0.52 0.155 0.52 0.155 0.06 0 0.06 0 -0.06 8.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 8.1 1.335 7.61 1.335 7.61 1.275 8.04 1.275 8.04 1.175 7.22 1.175 7.22 0.935 7.16 0.935 7.16 0.875 7.28 0.875 7.28 1.115 8.04 1.115 8.04 0.555 7.935 0.555 7.935 0.435 7.995 0.435 7.995 0.495 8.1 0.495 ;
      POLYGON 7.255 0.42 6.9 0.42 6.9 1.035 7.12 1.035 7.12 1.395 7.06 1.395 7.06 1.095 6.84 1.095 6.84 0.4 5.56 0.4 5.56 0.605 5.72 0.605 5.72 0.965 5.78 0.965 5.78 1.025 5.66 1.025 5.66 0.665 5.5 0.665 5.5 0.34 7.255 0.34 ;
      POLYGON 6.545 1.095 6.37 1.095 6.37 1.055 6.11 1.055 6.11 1.41 4.96 1.41 4.96 1.12 4.64 1.12 4.64 1.18 4.04 1.18 4.04 1.055 3.4 1.055 3.4 1.19 3.02 1.19 3.02 0.36 2.7 0.36 2.7 0.68 2.58 0.68 2.58 0.62 2.64 0.62 2.64 0.3 3.08 0.3 3.08 1.13 3.34 1.13 3.34 0.995 4.1 0.995 4.1 1.12 4.58 1.12 4.58 1.06 5.02 1.06 5.02 1.35 6.05 1.35 6.05 0.65 6.09 0.65 6.09 0.5 6.525 0.5 6.525 0.56 6.15 0.56 6.15 0.71 6.11 0.71 6.11 0.995 6.43 0.995 6.43 1.035 6.545 1.035 ;
      POLYGON 5.99 0.56 5.95 0.56 5.95 1.25 5.12 1.25 5.12 0.76 4.8 0.76 4.8 0.8 4.36 0.8 4.36 0.715 3.34 0.715 3.34 0.655 4.42 0.655 4.42 0.74 4.74 0.74 4.74 0.7 5.24 0.7 5.24 0.76 5.18 0.76 5.18 1.19 5.5 1.19 5.5 0.765 5.56 0.765 5.56 1.19 5.89 1.19 5.89 0.56 5.87 0.56 5.87 0.5 5.99 0.5 ;
      POLYGON 5.4 1.09 5.28 1.09 5.28 1.03 5.34 1.03 5.34 0.6 4.64 0.6 4.64 0.64 4.52 0.64 4.52 0.58 4.58 0.58 4.58 0.54 5.215 0.54 5.215 0.39 5.275 0.39 5.275 0.54 5.4 0.54 ;
      POLYGON 5.02 0.92 4.96 0.92 4.96 0.96 4.48 0.96 4.48 1.02 4.42 1.02 4.42 0.96 4.2 0.96 4.2 0.895 3.24 0.895 3.24 1.03 3.18 1.03 3.18 0.43 3.24 0.43 3.24 0.495 4.36 0.495 4.36 0.42 4.48 0.42 4.48 0.48 4.42 0.48 4.42 0.555 3.24 0.555 3.24 0.835 4.26 0.835 4.26 0.9 4.9 0.9 4.9 0.86 5.02 0.86 ;
      POLYGON 4.66 0.425 4.58 0.425 4.58 0.32 4.26 0.32 4.26 0.395 4.14 0.395 4.14 0.315 4.18 0.315 4.18 0.24 4.66 0.24 ;
      POLYGON 2.92 1.19 2.86 1.19 2.86 0.84 1.88 0.84 1.88 0.715 1.635 0.715 1.635 0.65 1.39 0.65 1.39 0.385 0.785 0.385 0.785 0.775 0.725 0.775 0.725 0.325 1.45 0.325 1.45 0.59 1.695 0.59 1.695 0.655 1.94 0.655 1.94 0.78 2.8 0.78 2.8 0.46 2.92 0.46 ;
      POLYGON 2.6 1.22 2.54 1.22 2.54 1.16 1.815 1.16 1.815 1.22 1.755 1.22 1.755 1.1 2.6 1.1 ;
      POLYGON 2.54 0.52 2.48 0.52 2.48 0.67 2.04 0.67 2.04 0.555 1.93 0.555 1.93 0.475 2.12 0.475 2.12 0.59 2.4 0.59 2.4 0.44 2.54 0.44 ;
      POLYGON 2.3 0.49 2.22 0.49 2.22 0.375 1.83 0.375 1.83 0.49 1.75 0.49 1.75 0.295 2.3 0.295 ;
      POLYGON 2.09 1.48 1.56 1.48 1.56 1.16 1.1 1.16 1.1 0.995 1.045 0.995 1.045 0.485 1.225 0.485 1.225 0.545 1.105 0.545 1.105 0.935 1.16 0.935 1.16 1.1 1.62 1.1 1.62 1.42 2.09 1.42 ;
      POLYGON 1.3 1.55 0.885 1.55 0.885 0.935 0.56 0.935 0.56 0.73 0.62 0.73 0.62 0.875 0.885 0.875 0.885 0.485 0.945 0.485 0.945 1.49 1.3 1.49 ;
  END
END SDFFSRHQX2

MACRO SDFFSRHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRHQX4 0 0 ;
  SIZE 8.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 18.381877 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.135 1.34 4.46 1.34 4.46 1.285 4.14 1.285 4.14 1.405 3.28 1.405 3.28 1.065 3.165 1.065 3.165 1.085 3.035 1.085 3.035 1.065 2.89 1.065 2.89 1.005 3.34 1.005 3.34 1.345 4.08 1.345 4.08 1.225 4.52 1.225 4.52 1.28 5.135 1.28 ;
    END
  END SN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.99669975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.4 0.745 8.32 0.745 8.32 0.705 7.46 0.705 7.46 0.625 8.4 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.135 0.965 7.715 0.965 7.715 0.835 7.835 0.835 7.835 0.805 8.135 0.805 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.98 1.085 6.86 1.085 6.86 0.625 6.94 0.625 6.94 0.865 6.98 0.865 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.76 1.07 6.68 1.07 6.68 0.895 6.435 0.895 6.435 0.815 6.76 0.815 ;
    END
  END CK
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.75 1.74 1.25 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.74565 LAYER Metal1 ;
    ANTENNADIFFAREA 5.21915 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.417375 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.3702305 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 88.43845475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.905 0.645 0.86 0.645 0.86 0.9 0.905 0.9 0.905 1.29 0.845 1.29 0.845 0.96 0.8 0.96 0.8 0.705 0.495 0.705 0.495 1.29 0.435 1.29 0.435 0.54 0.495 0.54 0.495 0.625 0.565 0.625 0.565 0.645 0.8 0.645 0.8 0.585 0.845 0.585 0.845 0.525 0.905 0.525 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.6 1.77 0 1.77 0 1.65 0.23 1.65 0.23 0.9 0.29 0.9 0.29 1.65 0.64 1.65 0.64 0.9 0.7 0.9 0.7 1.65 1.05 1.65 1.05 0.98 1.11 0.98 1.11 1.65 1.49 1.65 1.49 1.51 1.55 1.51 1.55 1.65 2.15 1.65 2.15 1.51 2.21 1.51 2.21 1.65 2.79 1.65 2.79 1.54 2.91 1.54 2.91 1.65 4.24 1.65 4.24 1.385 4.36 1.385 4.36 1.445 4.3 1.445 4.3 1.65 5.26 1.65 5.26 1.25 5.38 1.25 5.38 1.31 5.32 1.31 5.32 1.65 6.32 1.65 6.32 1.345 6.38 1.345 6.38 1.65 7.18 1.65 7.18 1.22 7.24 1.22 7.24 1.65 7.8 1.65 7.8 1.235 7.86 1.235 7.86 1.65 8.47 1.65 8.47 0.995 8.53 0.995 8.53 1.65 8.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.6 0.06 8.53 0.06 8.53 0.545 8.47 0.545 8.47 0.06 7.765 0.06 7.765 0.305 7.825 0.305 7.825 0.365 7.705 0.365 7.705 0.06 7.085 0.06 7.085 0.17 6.965 0.17 6.965 0.06 6.56 0.06 6.56 0.17 6.44 0.17 6.44 0.06 5.405 0.06 5.405 0.365 5.465 0.365 5.465 0.425 5.345 0.425 5.345 0.06 3.07 0.06 3.07 0.2 3.01 0.2 3.01 0.06 1.55 0.06 1.55 0.49 1.43 0.49 1.43 0.43 1.49 0.43 1.49 0.06 1.11 0.06 1.11 0.52 1.05 0.52 1.05 0.06 0.7 0.06 0.7 0.52 0.64 0.52 0.64 0.06 0.29 0.06 0.29 0.52 0.23 0.52 0.23 0.06 0 0.06 0 -0.06 8.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 8.355 1.085 8.295 1.085 8.295 1.125 7.555 1.125 7.555 0.865 7.3 0.865 7.3 0.685 7.24 0.685 7.24 0.625 7.3 0.625 7.3 0.465 8.29 0.465 8.29 0.525 7.36 0.525 7.36 0.805 7.615 0.805 7.615 1.065 8.235 1.065 8.235 1.025 8.355 1.025 ;
      POLYGON 7.55 1.345 7.49 1.345 7.49 1.285 7.395 1.285 7.395 1.025 7.08 1.025 7.08 0.365 5.95 0.365 5.95 0.455 5.945 0.455 5.945 1.18 5.885 1.18 5.885 0.305 7.425 0.305 7.425 0.365 7.14 0.365 7.14 0.965 7.455 0.965 7.455 1.225 7.55 1.225 ;
      POLYGON 7.065 1.245 6.22 1.245 6.22 1.37 5.505 1.37 5.505 1.15 4.62 1.15 4.62 1.125 3.98 1.125 3.98 1.245 3.6 1.245 3.6 0.425 3.28 0.425 3.28 0.745 3.16 0.745 3.16 0.685 3.22 0.685 3.22 0.365 3.66 0.365 3.66 1.185 3.92 1.185 3.92 1.065 4.68 1.065 4.68 1.09 5.505 1.09 5.505 0.93 5.625 0.93 5.625 0.99 5.565 0.99 5.565 1.31 6.16 1.31 6.16 1.185 6.275 1.185 6.275 0.745 6.225 0.745 6.225 0.625 6.28 0.625 6.28 0.465 6.715 0.465 6.715 0.525 6.34 0.525 6.34 0.685 6.335 0.685 6.335 1.185 7.065 1.185 ;
      POLYGON 6.18 0.525 6.115 0.525 6.115 0.96 6.175 0.96 6.175 1.02 6.055 1.02 6.055 0.86 6.045 0.86 6.045 0.74 6.055 0.74 6.055 0.465 6.18 0.465 ;
      POLYGON 5.785 1.15 5.74 1.15 5.74 1.21 5.68 1.21 5.68 1.09 5.725 1.09 5.725 0.67 5.1 0.67 5.1 0.61 5.685 0.61 5.685 0.42 5.785 0.42 ;
      POLYGON 5.625 0.83 4.94 0.83 4.94 0.795 3.92 0.795 3.92 0.735 5 0.735 5 0.77 5.625 0.77 ;
      POLYGON 5.405 0.99 4.78 0.99 4.78 0.965 3.82 0.965 3.82 1.085 3.76 1.085 3.76 0.495 3.82 0.495 3.82 0.575 4.765 0.575 4.765 0.5 4.885 0.5 4.885 0.56 4.825 0.56 4.825 0.635 3.82 0.635 3.82 0.905 4.84 0.905 4.84 0.93 5.405 0.93 ;
      POLYGON 5.065 0.505 4.985 0.505 4.985 0.4 4.665 0.4 4.665 0.475 4.545 0.475 4.545 0.395 4.585 0.395 4.585 0.32 5.065 0.32 ;
      POLYGON 3.5 1.245 3.44 1.245 3.44 0.905 2.79 0.905 2.79 1.06 2.15 1.06 2.15 1.41 1.415 1.41 1.415 0.82 1.475 0.82 1.475 1.35 2.09 1.35 2.09 1 2.73 1 2.73 0.845 3.38 0.845 3.38 0.525 3.5 0.525 ;
      POLYGON 3.18 1.28 2.585 1.28 2.585 1.16 2.665 1.16 2.665 1.2 3.06 1.2 3.06 1.185 3.18 1.185 ;
      POLYGON 3.18 1.55 3.01 1.55 3.01 1.44 2.31 1.44 2.31 1.38 3.07 1.38 3.07 1.49 3.18 1.49 ;
      POLYGON 3.12 0.585 2.85 0.585 2.85 0.42 2.53 0.42 2.53 0.495 2.41 0.495 2.41 0.435 2.47 0.435 2.47 0.36 2.91 0.36 2.91 0.525 3.12 0.525 ;
      POLYGON 2.75 0.655 2.63 0.655 2.63 0.9 2.09 0.9 2.09 0.58 2.03 0.58 2.03 0.52 2.15 0.52 2.15 0.84 2.57 0.84 2.57 0.595 2.63 0.595 2.63 0.52 2.75 0.52 ;
      POLYGON 2.47 0.74 2.25 0.74 2.25 0.415 1.71 0.415 1.71 0.65 1.315 0.65 1.315 1.29 1.255 1.29 1.255 0.8 0.96 0.8 0.96 0.74 1.255 0.74 1.255 0.485 1.315 0.485 1.315 0.59 1.65 0.59 1.65 0.355 2.31 0.355 2.31 0.68 2.47 0.68 ;
      POLYGON 1.99 0.845 1.92 0.845 1.92 1.1 1.84 1.1 1.84 0.595 1.81 0.595 1.81 0.515 1.93 0.515 1.93 0.595 1.92 0.595 1.92 0.765 1.99 0.765 ;
  END
END SDFFSRHQX4

MACRO SDFFSRHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRHQX8 0 0 ;
  SIZE 9.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.5148515 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.34 0.73 9.26 0.73 9.26 0.66 8.46 0.66 8.46 0.88 8.4 0.88 8.4 0.6 9.34 0.6 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.16 0.96 8.78 0.96 8.78 0.82 8.835 0.82 8.835 0.76 9.16 0.76 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 8.06 0.445 8.14 0.945 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.96 0.88 7.88 0.88 7.88 0.705 7.635 0.705 7.635 0.625 7.96 0.625 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 24.789644 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 1.34 5.24 1.34 5.24 1.195 4.92 1.195 4.92 1.365 4.06 1.365 4.06 1.015 3.12 1.015 3.12 0.92 3.06 0.92 3.06 0.79 3.14 0.79 3.14 0.815 3.18 0.815 3.18 0.955 4.12 0.955 4.12 1.305 4.86 1.305 4.86 1.135 5.3 1.135 5.3 1.28 6 1.28 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.96 0.87 2.765 0.87 2.765 0.975 2.565 0.975 2.565 0.79 2.96 0.79 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.439975 LAYER Metal1 ;
    ANTENNADIFFAREA 6.05495 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.574875 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.46288325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 74.5153295 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.37 0.65 1.325 0.65 1.325 0.9 1.37 0.9 1.37 1.345 1.31 1.345 1.31 0.96 1.265 0.96 1.265 0.8 0.96 0.8 0.96 1.345 0.9 1.345 0.9 0.66 0.55 0.66 0.55 1.345 0.49 1.345 0.49 0.66 0.14 0.66 0.14 1.345 0.08 1.345 0.08 0.73 0.06 0.73 0.06 0.6 0.08 0.6 0.08 0.54 0.14 0.54 0.14 0.6 0.49 0.6 0.49 0.54 0.55 0.54 0.55 0.6 0.9 0.6 0.9 0.54 0.96 0.54 0.96 0.74 1.265 0.74 1.265 0.59 1.31 0.59 1.31 0.53 1.37 0.53 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.6 1.77 0 1.77 0 1.65 0.285 1.65 0.285 0.9 0.345 0.9 0.345 1.65 0.695 1.65 0.695 0.9 0.755 0.9 0.755 1.65 1.105 1.65 1.105 0.9 1.165 0.9 1.165 1.65 1.515 1.65 1.515 0.955 1.575 0.955 1.575 1.65 1.925 1.65 1.925 1.045 1.985 1.045 1.985 1.65 2.855 1.65 2.855 1.295 2.975 1.295 2.975 1.355 2.915 1.355 2.915 1.65 3.67 1.65 3.67 1.275 3.79 1.275 3.79 1.335 3.73 1.335 3.73 1.65 5.08 1.65 5.08 1.355 5.02 1.355 5.02 1.295 5.14 1.295 5.14 1.65 6.1 1.65 6.1 1.22 6.22 1.22 6.22 1.28 6.16 1.28 6.16 1.65 7.57 1.65 7.57 1.14 7.63 1.14 7.63 1.65 8.06 1.65 8.06 1.045 8.12 1.045 8.12 1.65 8.835 1.65 8.835 1.22 8.895 1.22 8.895 1.65 9.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.6 0.06 9.01 0.06 9.01 0.5 8.95 0.5 8.95 0.06 8.21 0.06 8.21 0.17 8.09 0.17 8.09 0.06 7.545 0.06 7.545 0.17 7.425 0.17 7.425 0.06 6.215 0.06 6.215 0.425 6.155 0.425 6.155 0.06 3.04 0.06 3.04 0.53 2.92 0.53 2.92 0.47 2.98 0.47 2.98 0.06 1.985 0.06 1.985 0.485 1.925 0.485 1.925 0.06 1.575 0.06 1.575 0.485 1.515 0.485 1.515 0.06 1.165 0.06 1.165 0.485 1.105 0.485 1.105 0.06 0.755 0.06 0.755 0.485 0.695 0.485 0.695 0.06 0.345 0.06 0.345 0.485 0.285 0.485 0.285 0.06 0 0.06 0 -0.06 9.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 9.5 1.28 9.01 1.28 9.01 1.22 9.44 1.22 9.44 1.12 8.62 1.12 8.62 0.88 8.56 0.88 8.56 0.82 8.68 0.82 8.68 1.06 9.44 1.06 9.44 0.5 9.335 0.5 9.335 0.38 9.395 0.38 9.395 0.44 9.5 0.44 ;
      POLYGON 8.645 0.38 8.3 0.38 8.3 0.98 8.52 0.98 8.52 1.34 8.46 1.34 8.46 1.04 8.24 1.04 8.24 0.345 6.92 0.345 6.92 0.675 7.14 0.675 7.14 1.065 7.02 1.065 7.02 1.005 7.08 1.005 7.08 0.735 6.86 0.735 6.86 0.285 8.645 0.285 ;
      POLYGON 7.945 1.04 7.47 1.04 7.47 1.41 6.32 1.41 6.32 1.12 6 1.12 6 1.18 5.4 1.18 5.4 1.035 4.76 1.035 4.76 1.205 4.38 1.205 4.38 0.655 4.44 0.655 4.44 0.365 4.12 0.365 4.12 0.695 4 0.695 4 0.635 4.06 0.635 4.06 0.305 4.5 0.305 4.5 0.715 4.44 0.715 4.44 1.145 4.7 1.145 4.7 0.975 5.46 0.975 5.46 1.12 5.94 1.12 5.94 1.06 6.38 1.06 6.38 1.35 7.41 1.35 7.41 0.46 7.915 0.46 7.915 0.52 7.47 0.52 7.47 0.98 7.945 0.98 ;
      POLYGON 7.31 1.25 6.48 1.25 6.48 0.76 6.16 0.76 6.16 0.8 5.72 0.8 5.72 0.715 4.76 0.715 4.76 0.655 5.78 0.655 5.78 0.74 6.1 0.74 6.1 0.7 6.6 0.7 6.6 0.76 6.54 0.76 6.54 1.19 6.86 1.19 6.86 0.835 6.98 0.835 6.98 0.895 6.92 0.895 6.92 1.19 7.25 1.19 7.25 0.505 7.19 0.505 7.19 0.445 7.31 0.445 ;
      POLYGON 6.76 1.09 6.64 1.09 6.64 1.03 6.7 1.03 6.7 0.6 6 0.6 6 0.64 5.88 0.64 5.88 0.58 5.94 0.58 5.94 0.54 6.575 0.54 6.575 0.39 6.635 0.39 6.635 0.54 6.76 0.54 ;
      POLYGON 6.38 0.92 6.32 0.92 6.32 0.96 5.84 0.96 5.84 1.02 5.78 1.02 5.78 0.96 5.56 0.96 5.56 0.875 4.6 0.875 4.6 1.045 4.54 1.045 4.54 0.815 4.6 0.815 4.6 0.435 4.66 0.435 4.66 0.495 5.66 0.495 5.66 0.42 5.78 0.42 5.78 0.48 5.72 0.48 5.72 0.555 4.66 0.555 4.66 0.815 5.62 0.815 5.62 0.9 6.26 0.9 6.26 0.86 6.38 0.86 ;
      POLYGON 6.005 0.425 5.925 0.425 5.925 0.32 5.56 0.32 5.56 0.395 5.44 0.395 5.44 0.315 5.48 0.315 5.48 0.24 6.005 0.24 ;
      POLYGON 4.34 0.525 4.28 0.525 4.28 1.205 4.22 1.205 4.22 0.855 3.28 0.855 3.28 0.69 2.76 0.69 2.76 0.365 2.145 0.365 2.145 0.785 2.085 0.785 2.085 0.305 2.82 0.305 2.82 0.63 3.34 0.63 3.34 0.795 4.22 0.795 4.22 0.465 4.34 0.465 ;
      POLYGON 3.96 0.535 3.885 0.535 3.885 0.695 3.44 0.695 3.44 0.48 3.52 0.48 3.52 0.615 3.805 0.615 3.805 0.455 3.96 0.455 ;
      POLYGON 3.96 1.235 3.9 1.235 3.9 1.175 3.295 1.175 3.295 1.235 3.235 1.235 3.235 1.115 3.96 1.115 ;
      POLYGON 3.705 0.515 3.625 0.515 3.625 0.38 3.315 0.38 3.315 0.515 3.235 0.515 3.235 0.3 3.705 0.3 ;
      POLYGON 3.57 1.46 3.075 1.46 3.075 1.195 2.65 1.195 2.65 1.135 2.405 1.135 2.405 0.525 2.6 0.525 2.6 0.465 2.66 0.465 2.66 0.585 2.465 0.585 2.465 1.075 2.71 1.075 2.71 1.135 3.135 1.135 3.135 1.4 3.57 1.4 ;
      POLYGON 2.755 1.495 2.13 1.495 2.13 1.045 2.245 1.045 2.245 0.945 1.78 0.945 1.78 1.345 1.72 1.345 1.72 0.805 1.425 0.805 1.425 0.745 1.72 0.745 1.72 0.505 1.78 0.505 1.78 0.885 2.245 0.885 2.245 0.505 2.305 0.505 2.305 1.105 2.19 1.105 2.19 1.435 2.755 1.435 ;
  END
END SDFFSRHQX8

MACRO SDFFSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRX1 0 0 ;
  SIZE 7.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.965675 LAYER Metal1 ;
    ANTENNADIFFAREA 4.021075 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2691 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.736808 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 112.28539575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.955 0.485 0.94 0.485 0.94 0.83 0.955 0.83 0.955 1.43 0.895 1.43 0.895 0.89 0.88 0.89 0.88 0.73 0.86 0.73 0.86 0.6 0.88 0.6 0.88 0.44 0.895 0.44 0.895 0.365 0.955 0.365 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.965675 LAYER Metal1 ;
    ANTENNADIFFAREA 4.021075 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2691 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.736808 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 112.28539575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.32 1.29 0.24 1.29 0.24 0.73 0.06 0.73 0.06 0.6 0.24 0.6 0.24 0.54 0.32 0.54 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.14 0.745 7.08 0.745 7.08 0.715 6.415 0.715 6.415 1 6.355 1 6.355 0.655 6.675 0.655 6.675 0.595 6.735 0.595 6.735 0.655 6.835 0.655 6.835 0.625 7.14 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.98 0.93 6.515 0.93 6.515 0.85 6.635 0.85 6.635 0.815 6.98 0.815 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.595 0.815 6.095 0.895 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.095 1.075 5.765 1.075 5.765 1.085 5.605 1.085 5.605 1.005 5.685 1.005 5.685 0.995 6.095 0.995 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 27.45370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.375 3.885 1.375 3.885 1.215 2.985 1.215 2.985 0.985 2.035 0.985 2.035 0.875 1.995 0.875 1.995 0.815 2.165 0.815 2.165 0.925 3.045 0.925 3.045 1.155 3.945 1.155 3.945 1.315 4.4 1.315 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.71 1.34 1.21 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.4 1.77 0 1.77 0 1.65 0.465 1.65 0.465 0.995 0.525 0.995 0.525 1.65 1.1 1.65 1.1 1.31 1.16 1.31 1.16 1.65 1.865 1.65 1.865 1.51 1.925 1.51 1.925 1.65 2.505 1.65 2.505 1.425 2.625 1.425 2.625 1.485 2.565 1.485 2.565 1.65 3.495 1.65 3.495 1.54 3.615 1.54 3.615 1.65 4.5 1.65 4.5 1.51 4.56 1.51 4.56 1.65 5.35 1.65 5.35 1.54 5.47 1.54 5.47 1.65 5.935 1.65 5.935 1.285 6.055 1.285 6.055 1.345 5.995 1.345 5.995 1.65 6.845 1.65 6.845 1.255 6.905 1.255 6.905 1.65 7.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.4 0.06 6.98 0.06 6.98 0.495 6.92 0.495 6.92 0.06 6.23 0.06 6.23 0.395 6.11 0.395 6.11 0.335 6.17 0.335 6.17 0.06 5.47 0.06 5.47 0.17 5.35 0.17 5.35 0.06 4.49 0.06 4.49 0.575 4.43 0.575 4.43 0.06 1.955 0.06 1.955 0.17 1.835 0.17 1.835 0.06 1.16 0.06 1.16 0.45 1.1 0.45 1.1 0.06 0.525 0.06 0.525 0.635 0.465 0.635 0.465 0.06 0 0.06 0 -0.06 7.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.36 0.49 7.3 0.49 7.3 1.09 7.205 1.09 7.205 1.28 7.145 1.28 7.145 1.09 6.515 1.09 6.515 1.03 7.24 1.03 7.24 0.43 7.36 0.43 ;
      POLYGON 6.67 0.495 6.575 0.495 6.575 0.555 6.255 0.555 6.255 1.19 6.49 1.19 6.49 1.31 6.43 1.31 6.43 1.25 6.195 1.25 6.195 0.555 5.95 0.555 5.95 0.415 5.005 0.415 5.005 1.125 4.945 1.125 4.945 0.355 6.01 0.355 6.01 0.495 6.515 0.495 6.515 0.435 6.61 0.435 6.61 0.375 6.67 0.375 ;
      POLYGON 5.85 0.585 5.495 0.585 5.495 0.735 5.395 0.735 5.395 1.245 5.76 1.245 5.76 1.185 5.82 1.185 5.82 1.305 4.78 1.305 4.78 1.445 4.66 1.445 4.66 1.305 4.55 1.305 4.55 1.215 4.045 1.215 4.045 1.055 3.835 1.055 3.835 0.895 3.74 0.895 3.74 0.835 3.895 0.835 3.895 0.995 4.105 0.995 4.105 1.155 4.61 1.155 4.61 1.245 5.335 1.245 5.335 0.795 5.275 0.795 5.275 0.675 5.435 0.675 5.435 0.525 5.85 0.525 ;
      POLYGON 5.235 0.575 5.165 0.575 5.165 1.005 5.235 1.005 5.235 1.065 5.105 1.065 5.105 0.515 5.235 0.515 ;
      POLYGON 4.83 1.095 4.71 1.095 4.71 0.735 4.155 0.735 4.155 0.675 4.74 0.675 4.74 0.48 4.8 0.48 4.8 1.035 4.83 1.035 ;
      POLYGON 4.585 0.895 4.265 0.895 4.265 0.995 4.325 0.995 4.325 1.055 4.205 1.055 4.205 0.895 3.995 0.895 3.995 0.735 3.64 0.735 3.64 1.05 3.365 1.05 3.365 0.99 3.58 0.99 3.58 0.705 3.465 0.705 3.465 0.54 3.525 0.54 3.525 0.645 3.64 0.645 3.64 0.675 3.995 0.675 3.995 0.48 4.055 0.48 4.055 0.835 4.585 0.835 ;
      POLYGON 4.285 0.575 4.225 0.575 4.225 0.38 3.88 0.38 3.88 0.545 3.76 0.545 3.76 0.485 3.82 0.485 3.82 0.32 4.285 0.32 ;
      POLYGON 3.785 1.375 2.725 1.375 2.725 1.325 2.405 1.325 2.405 1.385 2.345 1.385 2.345 1.325 1.795 1.325 1.795 1.43 1.335 1.43 1.335 1.31 1.44 1.31 1.44 0.49 1.42 0.49 1.42 0.355 1.48 0.355 1.48 0.43 1.5 0.43 1.5 1.37 1.735 1.37 1.735 1.265 2.785 1.265 2.785 1.315 3.785 1.315 ;
      POLYGON 3.48 0.865 3.305 0.865 3.305 0.265 3.05 0.265 3.05 0.205 3.365 0.205 3.365 0.805 3.48 0.805 ;
      POLYGON 3.265 1.05 3.145 1.05 3.145 0.825 2.37 0.825 2.37 0.715 1.76 0.715 1.76 0.655 2.43 0.655 2.43 0.765 3.145 0.765 3.145 0.54 3.205 0.54 3.205 0.99 3.265 0.99 ;
      POLYGON 3.01 0.665 2.53 0.665 2.53 0.53 2.49 0.53 2.49 0.45 2.61 0.45 2.61 0.585 2.93 0.585 2.93 0.54 3.01 0.54 ;
      RECT 2.07 1.085 2.885 1.165 ;
      POLYGON 2.83 0.485 2.71 0.485 2.71 0.35 2.39 0.35 2.39 0.49 2.07 0.49 2.07 0.43 2.33 0.43 2.33 0.29 2.77 0.29 2.77 0.425 2.83 0.425 ;
      POLYGON 2.23 0.325 2.115 0.325 2.115 0.33 1.69 0.33 1.69 0.555 1.66 0.555 1.66 0.815 1.69 0.815 1.69 1.08 1.63 1.08 1.63 0.875 1.6 0.875 1.6 0.495 1.63 0.495 1.63 0.255 1.32 0.255 1.32 0.61 1.16 0.61 1.16 0.73 1.04 0.73 1.04 0.55 1.26 0.55 1.26 0.195 1.69 0.195 1.69 0.27 2.055 0.27 2.055 0.265 2.23 0.265 ;
      POLYGON 0.755 1.02 0.675 1.02 0.675 0.815 0.42 0.815 0.42 0.735 0.675 0.735 0.675 0.54 0.755 0.54 ;
  END
END SDFFSRX1

MACRO SDFFSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRX2 0 0 ;
  SIZE 9.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.96315 LAYER Metal1 ;
    ANTENNADIFFAREA 5.1663 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.334575 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.83419275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 114.270343 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.76 0.63 8.7 0.63 8.7 1.305 8.64 1.305 8.64 0.73 8.46 0.73 8.46 0.6 8.54 0.6 8.54 0.67 8.64 0.67 8.64 0.57 8.76 0.57 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.96315 LAYER Metal1 ;
    ANTENNADIFFAREA 5.1663 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.334575 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.83419275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 114.270343 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.2 1.305 8.12 1.305 8.12 1.11 8.06 1.11 8.06 0.98 8.12 0.98 8.12 0.54 8.2 0.54 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.86 1.085 7.635 1.085 7.635 0.73 7.715 0.73 7.715 0.95 7.86 0.95 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2142 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.611111 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 72.5925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.61 0.755 3.365 0.755 3.365 0.8 3.205 0.8 3.205 0.625 3.365 0.625 3.365 0.675 3.61 0.675 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.525 1.74 1.025 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 0.73 1.46 0.73 1.46 0.68 1.36 0.68 1.36 0.87 1.28 0.87 1.28 0.6 1.54 0.6 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.685 1.07 0.605 1.07 0.605 0.92 0.46 0.92 0.46 0.715 0.685 0.715 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 21.388889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.18 1.03 1.12 1.03 1.12 0.29 0.715 0.29 0.715 0.555 0.775 0.555 0.775 0.56 0.86 0.56 0.86 0.62 0.74 0.62 0.74 0.615 0.34 0.615 0.34 0.73 0.26 0.73 0.26 0.6 0.28 0.6 0.28 0.555 0.655 0.555 0.655 0.23 1.18 0.23 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.4 1.77 0 1.77 0 1.65 0.41 1.65 0.41 1.33 0.47 1.33 0.47 1.65 1.44 1.65 1.44 1.285 1.5 1.285 1.5 1.65 2.15 1.65 2.15 1.54 2.27 1.54 2.27 1.65 3.245 1.65 3.245 1.51 3.305 1.51 3.305 1.65 4.08 1.65 4.08 1.475 4.02 1.475 4.02 1.415 4.14 1.415 4.14 1.65 5.465 1.65 5.465 1.475 5.405 1.475 5.405 1.415 5.525 1.415 5.525 1.65 6.93 1.65 6.93 1.55 6.87 1.55 6.87 1.49 6.99 1.49 6.99 1.65 7.9 1.65 7.9 1.185 7.96 1.185 7.96 1.65 8.425 1.65 8.425 0.915 8.485 0.915 8.485 1.65 8.845 1.65 8.845 1.01 8.905 1.01 8.905 1.65 9.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.4 0.06 9.09 0.06 9.09 0.17 8.97 0.17 8.97 0.06 8.495 0.06 8.495 0.17 8.375 0.17 8.375 0.06 7.96 0.06 7.96 0.17 7.84 0.17 7.84 0.06 7.145 0.06 7.145 0.54 7.085 0.54 7.085 0.06 3.42 0.06 3.42 0.17 3.3 0.17 3.3 0.06 2.155 0.06 2.155 0.635 2.095 0.635 2.095 0.06 1.405 0.06 1.405 0.455 1.345 0.455 1.345 0.06 0.415 0.06 0.415 0.455 0.355 0.455 0.355 0.06 0 0.06 0 -0.06 9.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 9.325 0.63 9.135 0.63 9.135 1.035 9.075 1.035 9.075 0.79 8.8 0.79 8.8 0.73 9.075 0.73 9.075 0.57 9.325 0.57 ;
      POLYGON 9.25 0.44 8.36 0.44 8.36 0.83 8.3 0.83 8.3 0.44 8.02 0.44 8.02 0.83 7.96 0.83 7.96 0.44 7.375 0.44 7.375 1.025 7.31 1.025 7.31 1.245 7.25 1.245 7.25 0.965 7.315 0.965 7.315 0.705 6.805 0.705 6.805 0.645 7.315 0.645 7.315 0.38 9.13 0.38 9.13 0.375 9.25 0.375 ;
      POLYGON 7.785 0.63 7.535 0.63 7.535 1.185 7.755 1.185 7.755 1.405 7.09 1.405 7.09 1.185 5.785 1.185 5.785 1.155 5.3 1.155 5.3 1.095 5.845 1.095 5.845 1.125 7.15 1.125 7.15 1.345 7.695 1.345 7.695 1.245 7.475 1.245 7.475 0.57 7.785 0.57 ;
      POLYGON 7.215 0.865 6.105 0.865 6.105 0.835 4.94 0.835 4.94 1.02 4.88 1.02 4.88 0.45 4.94 0.45 4.94 0.775 6.165 0.775 6.165 0.805 7.215 0.805 ;
      POLYGON 6.945 0.54 6.865 0.54 6.865 0.375 6.545 0.375 6.545 0.51 6.425 0.51 6.425 0.43 6.465 0.43 6.465 0.295 6.945 0.295 ;
      POLYGON 6.77 1.345 5.625 1.345 5.625 1.315 4.94 1.315 4.94 1.34 4.24 1.34 4.24 1.315 3.92 1.315 3.92 1.44 3.405 1.44 3.405 1.38 3.86 1.38 3.86 1.255 4.3 1.255 4.3 1.28 4.88 1.28 4.88 1.255 5.685 1.255 5.685 1.285 6.77 1.285 ;
      POLYGON 6.765 0.535 6.705 0.535 6.705 0.67 6.265 0.67 6.265 0.54 5.055 0.54 5.055 0.48 6.325 0.48 6.325 0.61 6.645 0.61 6.645 0.475 6.765 0.475 ;
      POLYGON 6.74 1.025 5.945 1.025 5.945 0.995 5.145 0.995 5.145 1.055 5.085 1.055 5.085 0.935 6.005 0.935 6.005 0.965 6.74 0.965 ;
      POLYGON 5.02 0.22 4.78 0.22 4.78 1.18 4.4 1.18 4.4 1.155 3.76 1.155 3.76 1.28 3.32 1.28 3.32 1.12 3.045 1.12 3.045 0.765 3.105 0.765 3.105 1.06 3.38 1.06 3.38 1.22 3.7 1.22 3.7 1.095 4.46 1.095 4.46 1.12 4.72 1.12 4.72 0.16 5.02 0.16 ;
      POLYGON 4.62 1.02 4.56 1.02 4.56 0.96 3.6 0.96 3.6 1.12 3.48 1.12 3.48 1.06 3.54 1.06 3.54 0.96 3.205 0.96 3.205 0.9 4.105 0.9 4.105 0.46 4.165 0.46 4.165 0.9 4.56 0.9 4.56 0.45 4.62 0.45 ;
      POLYGON 4.37 0.555 4.31 0.555 4.31 0.36 4.005 0.36 4.005 0.525 3.87 0.525 3.87 0.465 3.945 0.465 3.945 0.3 4.37 0.3 ;
      POLYGON 3.94 0.735 3.71 0.735 3.71 0.525 2.945 0.525 2.945 1.175 2.885 1.175 2.885 0.465 3.77 0.465 3.77 0.675 3.94 0.675 ;
      POLYGON 3.845 0.29 3.785 0.29 3.785 0.33 2.785 0.33 2.785 1 2.725 1 2.725 0.33 2.425 0.33 2.425 0.58 2.465 0.58 2.465 0.96 2.405 0.96 2.405 1.02 2.345 1.02 2.345 0.9 2.405 0.9 2.405 0.64 2.365 0.64 2.365 0.27 3.725 0.27 3.725 0.23 3.845 0.23 ;
      POLYGON 2.71 1.44 1.6 1.44 1.6 1.185 1.34 1.185 1.34 1.19 1.02 1.19 1.02 1.355 0.96 1.355 0.96 0.45 0.815 0.45 0.815 0.39 1.02 0.39 1.02 1.13 1.28 1.13 1.28 1.125 1.66 1.125 1.66 1.38 2.565 1.38 2.565 0.46 2.625 0.46 2.625 1.15 2.71 1.15 ;
      POLYGON 2.305 0.8 1.9 0.8 1.9 1.28 1.76 1.28 1.76 1.22 1.84 1.22 1.84 0.425 1.705 0.425 1.705 0.365 1.9 0.365 1.9 0.74 2.305 0.74 ;
      POLYGON 0.86 1.23 0.265 1.23 0.265 1.355 0.205 1.355 0.205 1.23 0.1 1.23 0.1 0.43 0.12 0.43 0.12 0.36 0.18 0.36 0.18 0.48 0.16 0.48 0.16 1.17 0.8 1.17 0.8 0.795 0.86 0.795 ;
  END
END SDFFSRX2

MACRO SDFFSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRX4 0 0 ;
  SIZE 9.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4135 LAYER Metal1 ;
    ANTENNADIFFAREA 5.55505 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4878 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.097786 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 87.109471 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.855 0.51 8.385 0.51 8.385 0.79 8.54 0.79 8.54 0.86 8.7 0.86 8.7 0.955 8.745 0.955 8.745 1.305 8.685 1.305 8.685 1.015 8.64 1.015 8.64 0.92 8.38 0.92 8.38 0.975 8.335 0.975 8.335 1.305 8.275 1.305 8.275 0.915 8.32 0.915 8.32 0.51 8.265 0.51 8.265 0.45 8.855 0.45 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4135 LAYER Metal1 ;
    ANTENNADIFFAREA 5.55505 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4878 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.097786 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 87.109471 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.915 0.51 7.54 0.51 7.54 0.915 7.885 0.915 7.885 1.305 7.825 1.305 7.825 0.975 7.475 0.975 7.475 1.305 7.415 1.305 7.415 0.915 7.46 0.915 7.46 0.79 7.48 0.79 7.48 0.51 7.325 0.51 7.325 0.45 7.915 0.45 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.815 0.895 4.575 0.895 4.575 0.555 4.655 0.555 4.655 0.815 4.815 0.815 ;
    END
  END RN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.475 0.895 4.235 0.895 4.235 0.815 4.31 0.815 4.31 0.555 4.39 0.555 4.39 0.815 4.475 0.815 ;
    END
  END SN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.765 0.705 1.535 0.705 1.535 0.895 1.455 0.895 1.455 0.625 1.765 0.625 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 1.01 1.26 1.01 1.26 0.805 1.185 0.805 1.185 0.585 1.265 0.585 1.265 0.725 1.34 0.725 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.605 0.98 0.2 0.98 0.2 0.805 0.365 0.805 0.365 0.9 0.605 0.9 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 19.25925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.145 0.965 1.025 0.965 1.025 0.32 0.68 0.32 0.68 0.625 0.765 0.625 0.765 0.705 0.62 0.705 0.62 0.645 0.36 0.645 0.36 0.705 0.3 0.705 0.3 0.585 0.62 0.585 0.62 0.26 1.085 0.26 1.085 0.905 1.145 0.905 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.6 1.77 0 1.77 0 1.65 0.43 1.65 0.43 1.24 0.49 1.24 0.49 1.65 1.295 1.65 1.295 1.27 1.415 1.27 1.415 1.33 1.355 1.33 1.355 1.65 2.82 1.65 2.82 1.54 2.94 1.54 2.94 1.65 3.305 1.65 3.305 1.54 3.425 1.54 3.425 1.65 4.435 1.65 4.435 1.375 4.375 1.375 4.375 1.315 4.495 1.315 4.495 1.65 6.145 1.65 6.145 1.185 6.205 1.185 6.205 1.65 6.66 1.65 6.66 1.185 6.72 1.185 6.72 1.65 7.07 1.65 7.07 0.995 7.13 0.995 7.13 1.65 7.62 1.65 7.62 1.075 7.68 1.075 7.68 1.65 8.03 1.65 8.03 0.915 8.09 0.915 8.09 1.65 8.48 1.65 8.48 1.02 8.54 1.02 8.54 1.65 8.89 1.65 8.89 0.96 8.95 0.96 8.95 1.65 9.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.6 0.06 9.235 0.06 9.235 0.37 9.115 0.37 9.115 0.31 9.175 0.31 9.175 0.06 8.62 0.06 8.62 0.17 8.5 0.17 8.5 0.06 8.15 0.06 8.15 0.17 8.03 0.17 8.03 0.06 7.68 0.06 7.68 0.17 7.56 0.17 7.56 0.06 7.005 0.06 7.005 0.365 7.065 0.365 7.065 0.425 6.945 0.425 6.945 0.06 6.625 0.06 6.625 0.455 6.565 0.455 6.565 0.06 4.51 0.06 4.51 0.235 4.57 0.235 4.57 0.295 4.45 0.295 4.45 0.06 2.99 0.06 2.99 0.17 2.87 0.17 2.87 0.06 1.31 0.06 1.31 0.485 1.25 0.485 1.25 0.06 0.49 0.06 0.49 0.485 0.43 0.485 0.43 0.06 0 0.06 0 -0.06 9.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 9.41 0.86 9.155 0.86 9.155 1.305 9.095 1.305 9.095 0.86 8.8 0.86 8.8 0.785 8.92 0.785 8.92 0.8 9.35 0.8 9.35 0.42 9.41 0.42 ;
      POLYGON 9.09 0.7 9.03 0.7 9.03 0.64 8.955 0.64 8.955 0.35 7.225 0.35 7.225 0.645 6.925 0.645 6.925 0.755 7.305 0.755 7.305 0.815 6.925 0.815 6.925 1.305 6.865 1.305 6.865 0.645 6.295 0.645 6.295 0.585 6.77 0.585 6.77 0.42 6.83 0.42 6.83 0.585 7.165 0.585 7.165 0.29 9.015 0.29 9.015 0.58 9.09 0.58 ;
      POLYGON 6.765 0.925 5.455 0.925 5.455 1.13 5.395 1.13 5.395 0.51 5.455 0.51 5.455 0.865 6.705 0.865 6.705 0.805 6.765 0.805 ;
      POLYGON 6.545 1.18 6.425 1.18 6.425 1.085 5.57 1.085 5.57 1.025 6.485 1.025 6.485 1.12 6.545 1.12 ;
      POLYGON 6.42 0.455 6.36 0.455 6.36 0.26 6.015 0.26 6.015 0.425 5.895 0.425 5.895 0.365 5.955 0.365 5.955 0.2 6.42 0.2 ;
      POLYGON 6.195 0.605 5.715 0.605 5.715 0.485 5.795 0.485 5.795 0.525 6.115 0.525 6.115 0.36 6.195 0.36 ;
      POLYGON 6.095 0.765 5.555 0.765 5.555 0.295 4.775 0.295 4.775 0.395 4.975 0.395 4.975 1.02 4.915 1.02 4.915 0.455 4.29 0.455 4.29 0.26 3.855 0.26 3.855 0.2 4.35 0.2 4.35 0.395 4.715 0.395 4.715 0.235 5.615 0.235 5.615 0.705 6.095 0.705 ;
      POLYGON 5.55 1.385 4.595 1.385 4.595 1.215 3.855 1.215 3.855 1.065 3.105 1.065 3.105 1.005 3.165 1.005 3.165 0.685 2.645 0.685 2.645 0.83 2.585 0.83 2.585 0.625 3.105 0.625 3.105 0.57 3.225 0.57 3.225 1.005 3.915 1.005 3.915 1.155 4.655 1.155 4.655 1.325 5.235 1.325 5.235 0.71 5.295 0.71 5.295 1.325 5.55 1.325 ;
      POLYGON 5.22 0.61 5.135 0.61 5.135 1.225 5.075 1.225 5.075 1.18 4.755 1.18 4.755 1.055 4.015 1.055 4.015 0.905 3.375 0.905 3.375 0.445 2.65 0.445 2.65 0.385 3.375 0.385 3.375 0.2 3.755 0.2 3.755 0.365 4.015 0.365 4.015 0.425 3.695 0.425 3.695 0.26 3.435 0.26 3.435 0.845 4.135 0.845 4.135 0.995 4.815 0.995 4.815 1.12 5.075 1.12 5.075 0.55 5.16 0.55 5.16 0.49 5.22 0.49 ;
      POLYGON 4.275 1.48 3.695 1.48 3.695 1.225 2.945 1.225 2.945 0.99 2.425 0.99 2.425 0.365 1.59 0.365 1.59 0.465 1.925 0.465 1.925 1.235 1.675 1.235 1.675 1.175 1.865 1.175 1.865 0.525 1.53 0.525 1.53 0.305 2.485 0.305 2.485 0.93 2.945 0.93 2.945 0.785 3.065 0.785 3.065 0.905 3.005 0.905 3.005 1.165 3.755 1.165 3.755 1.42 4.275 1.42 ;
      POLYGON 4.19 0.585 3.535 0.585 3.535 0.36 3.595 0.36 3.595 0.525 4.13 0.525 4.13 0.36 4.19 0.36 ;
      POLYGON 3.595 1.385 2.51 1.385 2.51 1.15 2.265 1.15 2.265 0.54 2.325 0.54 2.325 1.09 2.57 1.09 2.57 1.325 3.595 1.325 ;
      POLYGON 2.165 1.395 1.515 1.395 1.515 1.17 0.925 1.17 0.925 1.265 0.865 1.265 0.865 0.48 0.78 0.48 0.78 0.42 0.925 0.42 0.925 1.11 1.575 1.11 1.575 1.335 2.105 1.335 2.105 0.63 2.03 0.63 2.03 0.57 2.165 0.57 ;
      POLYGON 0.765 1.14 0.285 1.14 0.285 1.265 0.225 1.265 0.225 1.14 0.04 1.14 0.04 0.425 0.225 0.425 0.225 0.365 0.285 0.365 0.285 0.485 0.1 0.485 0.1 1.08 0.705 1.08 0.705 0.985 0.765 0.985 ;
  END
END SDFFSRX4

MACRO SDFFSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSRXL 0 0 ;
  SIZE 7.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9773 LAYER Metal1 ;
    ANTENNADIFFAREA 4.0338 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.243 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.36748975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 125.462963 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.995 0.635 0.94 0.635 0.94 1.255 0.88 1.255 0.88 0.73 0.86 0.73 0.86 0.6 0.88 0.6 0.88 0.55 0.935 0.55 0.935 0.515 0.995 0.515 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.028975 LAYER Metal1 ;
    ANTENNADIFFAREA 4.0338 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.243 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.580144 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 126.54321 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.31 0.62 0.26 0.62 0.26 0.9 0.31 0.9 0.31 1.02 0.23 1.02 0.23 0.99 0.18 0.99 0.18 0.73 0.06 0.73 0.06 0.6 0.16 0.6 0.16 0.53 0.23 0.53 0.23 0.405 0.31 0.405 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.324074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.365 0.715 6.775 0.715 6.775 1 6.715 1 6.715 0.655 6.895 0.655 6.895 0.595 6.955 0.595 6.955 0.655 7.235 0.655 7.235 0.625 7.275 0.625 7.275 0.595 7.335 0.595 7.335 0.625 7.365 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.035 0.815 7.275 0.985 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.455 1.175 6.375 1.175 6.375 0.895 6.235 0.895 6.235 0.815 6.455 0.815 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.775 1.005 6.275 1.085 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 27.5 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.485 1.4 4 1.4 4 1.24 3.09 1.24 3.09 1.01 2.305 1.01 2.305 0.895 2.1 0.895 2.1 0.835 2.235 0.835 2.235 0.815 2.365 0.815 2.365 0.95 3.15 0.95 3.15 1.18 4.06 1.18 4.06 1.34 4.485 1.34 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.39 1.13 1.245 1.13 1.245 1.085 1.04 1.085 1.04 0.9 1.365 0.9 1.365 0.995 1.39 0.995 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.6 1.77 0 1.77 0 1.65 0.455 1.65 0.455 0.995 0.515 0.995 0.515 1.65 1.145 1.65 1.145 1.23 1.205 1.23 1.205 1.65 1.97 1.65 1.97 1.51 2.03 1.51 2.03 1.65 2.61 1.65 2.61 1.49 2.73 1.49 2.73 1.55 2.67 1.55 2.67 1.65 3.61 1.65 3.61 1.54 3.73 1.54 3.73 1.65 4.585 1.65 4.585 1.51 4.645 1.51 4.645 1.65 5.585 1.65 5.585 1.345 5.705 1.345 5.705 1.405 5.645 1.405 5.645 1.65 6.3 1.65 6.3 1.275 6.42 1.275 6.42 1.335 6.36 1.335 6.36 1.65 7.14 1.65 7.14 1.245 7.2 1.245 7.2 1.65 7.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.6 0.06 7.2 0.06 7.2 0.52 7.14 0.52 7.14 0.06 6.39 0.06 6.39 0.395 6.27 0.395 6.27 0.335 6.33 0.335 6.33 0.06 5.64 0.06 5.64 0.17 5.52 0.17 5.52 0.06 4.615 0.06 4.615 0.6 4.555 0.6 4.555 0.06 2.06 0.06 2.06 0.17 1.94 0.17 1.94 0.06 1.205 0.06 1.205 0.635 1.145 0.635 1.145 0.06 0.545 0.06 0.545 0.2 0.485 0.2 0.485 0.06 0 0.06 0 -0.06 7.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.525 1.145 7.405 1.145 7.405 1.27 7.345 1.27 7.345 1.145 6.875 1.145 6.875 0.98 6.935 0.98 6.935 1.085 7.465 1.085 7.465 0.495 7.315 0.495 7.315 0.435 7.525 0.435 ;
      POLYGON 6.92 0.495 6.795 0.495 6.795 0.555 6.615 0.555 6.615 1.245 6.85 1.245 6.85 1.365 6.79 1.365 6.79 1.305 6.555 1.305 6.555 0.555 6.11 0.555 6.11 0.42 5.175 0.42 5.175 1.065 5.19 1.065 5.19 1.185 5.13 1.185 5.13 1.125 5.115 1.125 5.115 0.36 6.17 0.36 6.17 0.495 6.735 0.495 6.735 0.435 6.92 0.435 ;
      POLYGON 6.185 1.305 6.125 1.305 6.125 1.245 5.485 1.245 5.485 1.41 4.95 1.41 4.95 1.485 4.83 1.485 4.83 1.41 4.585 1.41 4.585 1.24 4.16 1.24 4.16 1.08 3.905 1.08 3.905 0.92 3.845 0.92 3.845 0.86 3.965 0.86 3.965 1.02 4.22 1.02 4.22 1.18 4.645 1.18 4.645 1.35 5.425 1.35 5.425 1.185 5.615 1.185 5.615 0.76 5.515 0.76 5.515 0.82 5.455 0.82 5.455 0.7 5.615 0.7 5.615 0.55 6.01 0.55 6.01 0.61 5.675 0.61 5.675 1.185 6.185 1.185 ;
      POLYGON 5.47 1.045 5.29 1.045 5.29 0.965 5.275 0.965 5.275 0.52 5.405 0.52 5.405 0.6 5.355 0.6 5.355 0.885 5.37 0.885 5.37 0.965 5.47 0.965 ;
      POLYGON 5.015 1.12 4.895 1.12 4.895 0.76 4.28 0.76 4.28 0.7 4.895 0.7 4.895 0.505 4.955 0.505 4.955 1.06 5.015 1.06 ;
      POLYGON 4.74 0.92 4.38 0.92 4.38 1.02 4.44 1.02 4.44 1.08 4.32 1.08 4.32 0.92 4.12 0.92 4.12 0.73 3.745 0.73 3.745 1.075 3.48 1.075 3.48 1.015 3.685 1.015 3.685 0.73 3.57 0.73 3.57 0.54 3.63 0.54 3.63 0.67 4.12 0.67 4.12 0.505 4.18 0.505 4.18 0.86 4.74 0.86 ;
      POLYGON 4.41 0.6 4.35 0.6 4.35 0.405 4.02 0.405 4.02 0.57 3.885 0.57 3.885 0.51 3.96 0.51 3.96 0.345 4.41 0.345 ;
      POLYGON 3.9 1.4 2.83 1.4 2.83 1.35 2.51 1.35 2.51 1.41 2.45 1.41 2.45 1.35 1.35 1.35 1.35 1.23 1.49 1.23 1.49 0.54 1.55 0.54 1.55 1.29 2.89 1.29 2.89 1.34 3.9 1.34 ;
      POLYGON 3.585 0.89 3.41 0.89 3.41 0.29 3.155 0.29 3.155 0.23 3.47 0.23 3.47 0.83 3.585 0.83 ;
      POLYGON 3.38 1.075 3.25 1.075 3.25 0.85 2.475 0.85 2.475 0.715 1.835 0.715 1.835 0.655 2.535 0.655 2.535 0.79 3.25 0.79 3.25 0.54 3.31 0.54 3.31 1.015 3.38 1.015 ;
      POLYGON 3.115 0.69 2.635 0.69 2.635 0.555 2.595 0.555 2.595 0.475 2.715 0.475 2.715 0.61 3.035 0.61 3.035 0.54 3.115 0.54 ;
      RECT 2.175 1.11 2.99 1.19 ;
      POLYGON 2.935 0.51 2.815 0.51 2.815 0.375 2.495 0.375 2.495 0.51 2.175 0.51 2.175 0.45 2.435 0.45 2.435 0.315 2.875 0.315 2.875 0.45 2.935 0.45 ;
      POLYGON 2.335 0.35 1.795 0.35 1.795 0.555 1.735 0.555 1.735 0.815 1.795 0.815 1.795 1.105 1.735 1.105 1.735 0.875 1.675 0.875 1.675 0.495 1.735 0.495 1.735 0.35 1.39 0.35 1.39 0.8 1.04 0.8 1.04 0.74 1.33 0.74 1.33 0.29 2.335 0.29 ;
      POLYGON 0.72 1.02 0.64 1.02 0.64 0.8 0.36 0.8 0.36 0.72 0.64 0.72 0.64 0.38 0.72 0.38 ;
  END
END SDFFSRXL

MACRO SDFFSX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSX1 0 0 ;
  SIZE 7 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.512 LAYER Metal1 ;
    ANTENNADIFFAREA 3.742225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2367 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.83734675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 113.25728775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.255 1.04 1.14 1.04 1.14 1.29 1.08 1.29 1.08 1.11 1.06 1.11 1.06 0.98 1.08 0.98 1.08 0.9 1.195 0.9 1.195 0.54 1.255 0.54 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.512 LAYER Metal1 ;
    ANTENNADIFFAREA 3.742225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2367 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.83734675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 113.25728775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 0.98 0.5 0.98 0.5 1.29 0.42 1.29 0.42 0.9 0.46 0.9 0.46 0.65 0.39 0.65 0.39 0.57 0.54 0.57 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.324074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.725 0.705 6.495 0.705 6.495 0.715 6.135 0.715 6.135 0.93 6.015 0.93 6.015 0.87 6.075 0.87 6.075 0.655 6.355 0.655 6.355 0.585 6.415 0.585 6.415 0.625 6.565 0.625 6.565 0.645 6.665 0.645 6.665 0.585 6.725 0.585 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.695 0.935 6.46 0.935 6.46 0.895 6.235 0.895 6.235 0.815 6.695 0.815 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.755 0.8 5.46 0.8 5.46 0.515 5.54 0.515 5.54 0.72 5.755 0.72 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.36 0.995 5.28 0.995 5.28 0.73 5.26 0.73 5.26 0.55 5.28 0.55 5.28 0.515 5.36 0.515 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 21.712963 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.515 0.39 3.455 0.39 3.455 0.41 3.015 0.41 3.015 0.385 2.295 0.385 2.295 0.815 2.365 0.815 2.365 0.895 1.855 0.895 1.855 0.835 2.235 0.835 2.235 0.325 3.075 0.325 3.075 0.35 3.395 0.35 3.395 0.33 3.515 0.33 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7 1.77 0 1.77 0 1.65 0.215 1.65 0.215 0.91 0.275 0.91 0.275 1.65 0.875 1.65 0.875 0.9 0.935 0.9 0.935 1.65 1.755 1.65 1.755 1.305 1.815 1.305 1.815 1.65 2.15 1.65 2.15 1.335 2.27 1.335 2.27 1.395 2.21 1.395 2.21 1.65 3.51 1.65 3.51 1.54 3.63 1.54 3.63 1.65 4.07 1.65 4.07 1.51 4.13 1.51 4.13 1.65 5.705 1.65 5.705 1.255 5.765 1.255 5.765 1.65 6.535 1.65 6.535 1.255 6.595 1.255 6.595 1.65 7 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7 0.06 6.65 0.06 6.65 0.415 6.59 0.415 6.59 0.06 5.52 0.06 5.52 0.415 5.46 0.415 5.46 0.06 4.155 0.06 4.155 0.375 4.095 0.375 4.095 0.06 3.295 0.06 3.295 0.25 3.175 0.25 3.175 0.19 3.235 0.19 3.235 0.06 1.87 0.06 1.87 0.57 1.81 0.57 1.81 0.06 0.935 0.06 0.935 0.52 0.875 0.52 0.875 0.06 0.245 0.06 0.245 0.2 0.185 0.2 0.185 0.06 0 0.06 0 -0.06 7 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.885 1.095 6.8 1.095 6.8 1.28 6.74 1.28 6.74 1.095 6.3 1.095 6.3 1.09 6.185 1.09 6.185 1.03 6.36 1.03 6.36 1.035 6.825 1.035 6.825 0.32 6.885 0.32 ;
      POLYGON 6.34 0.44 5.975 0.44 5.975 0.575 5.915 0.575 5.915 1.095 6.085 1.095 6.085 1.19 6.18 1.19 6.18 1.31 6.12 1.31 6.12 1.25 6.025 1.25 6.025 1.155 4.87 1.155 4.87 1.06 4.93 1.06 4.93 0.525 4.87 0.525 4.87 0.465 4.99 0.465 4.99 1.095 5.855 1.095 5.855 0.515 5.915 0.515 5.915 0.38 6.28 0.38 6.28 0.32 6.34 0.32 ;
      POLYGON 5.59 1.345 4.45 1.345 4.45 1.37 4.33 1.37 4.33 1.345 3.35 1.345 3.35 1.285 4.71 1.285 4.71 0.295 5.285 0.295 5.285 0.415 5.225 0.415 5.225 0.355 4.77 0.355 4.77 1.285 5.59 1.285 ;
      POLYGON 4.61 0.855 4.495 0.855 4.495 1.055 4.435 1.055 4.435 0.855 3.935 0.855 3.935 0.795 4.55 0.795 4.55 0.435 4.61 0.435 ;
      POLYGON 4.45 0.695 4.33 0.695 4.33 0.535 3.935 0.535 3.935 0.385 3.675 0.385 3.675 0.55 3.615 0.55 3.615 0.735 3.395 0.735 3.395 1.025 3.275 1.025 3.275 0.965 3.335 0.965 3.335 0.735 2.785 0.735 2.785 0.675 2.855 0.675 2.855 0.485 2.915 0.485 2.915 0.675 3.555 0.675 3.555 0.49 3.615 0.49 3.615 0.325 3.995 0.325 3.995 0.475 4.39 0.475 4.39 0.635 4.45 0.635 ;
      POLYGON 4.23 0.695 3.835 0.695 3.835 1.075 3.81 1.075 3.81 1.185 2.875 1.185 2.875 0.895 2.625 0.895 2.625 0.505 2.745 0.505 2.745 0.565 2.685 0.565 2.685 0.835 2.935 0.835 2.935 1.125 3.75 1.125 3.75 1.015 3.775 1.015 3.775 0.485 3.835 0.485 3.835 0.635 4.23 0.635 ;
      POLYGON 2.73 1.15 2.67 1.15 2.67 1.055 1.685 1.055 1.685 0.995 2.465 0.995 2.465 0.565 2.405 0.565 2.405 0.505 2.525 0.505 2.525 0.995 2.73 0.995 ;
      POLYGON 2.555 1.235 2.05 1.235 2.05 1.3 1.93 1.3 1.93 1.22 1.97 1.22 1.97 1.155 2.555 1.155 ;
      POLYGON 2.135 0.735 1.585 0.735 1.585 1.3 1.465 1.3 1.465 1.24 1.525 1.24 1.525 0.515 1.605 0.515 1.605 0.415 1.095 0.415 1.095 0.79 0.91 0.79 0.91 0.73 1.035 0.73 1.035 0.355 1.665 0.355 1.665 0.575 1.585 0.575 1.585 0.675 2.135 0.675 ;
      POLYGON 0.7 1.02 0.64 1.02 0.64 0.47 0.29 0.47 0.29 0.75 0.36 0.75 0.36 0.81 0.23 0.81 0.23 0.41 0.7 0.41 ;
  END
END SDFFSX1

MACRO SDFFSX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSX2 0 0 ;
  SIZE 6.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.51845 LAYER Metal1 ;
    ANTENNADIFFAREA 3.7621 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.302175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.6437495 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 89.7890295 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.145 1.29 1.065 1.29 1.065 0.73 1.06 0.73 1.06 0.6 1.065 0.6 1.065 0.54 1.145 0.54 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.47085 LAYER Metal1 ;
    ANTENNADIFFAREA 3.7621 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.302175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.48622475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 88.96500375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.34 1.29 0.28 1.29 0.28 0.73 0.26 0.73 0.26 0.6 0.28 0.6 0.28 0.54 0.34 0.54 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.87962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.505 0.685 6.365 0.685 6.365 0.705 5.95 0.705 5.95 1.085 5.83 1.085 5.83 1.025 5.89 1.025 5.89 0.645 6.105 0.645 6.105 0.585 6.165 0.585 6.165 0.625 6.505 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.61 1.055 6.27 1.055 6.27 0.975 6.435 0.975 6.435 0.815 6.61 0.815 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.63 0.63 5.54 0.63 5.54 0.765 5.46 0.765 5.46 0.63 5.265 0.63 5.265 0.55 5.63 0.55 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.165 1.085 5.035 1.085 5.035 1.005 5.045 1.005 5.045 0.635 5.165 0.635 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 24.39814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.505 0.39 3.445 0.39 3.445 0.55 3.005 0.55 3.005 0.375 2.295 0.375 2.295 0.815 2.365 0.815 2.365 0.895 1.855 0.895 1.855 0.835 2.235 0.835 2.235 0.315 3.065 0.315 3.065 0.49 3.385 0.49 3.385 0.33 3.505 0.33 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.8 1.77 0 1.77 0 1.65 0.075 1.65 0.075 0.9 0.135 0.9 0.135 1.65 0.485 1.65 0.485 1.17 0.545 1.17 0.545 1.65 0.85 1.65 0.85 1.285 0.91 1.285 0.91 1.65 1.32 1.65 1.32 1.51 1.38 1.51 1.38 1.65 1.71 1.65 1.71 1.305 1.77 1.305 1.77 1.65 2.105 1.65 2.105 1.335 2.225 1.335 2.225 1.395 2.165 1.395 2.165 1.65 3.5 1.65 3.5 1.54 3.62 1.54 3.62 1.65 4.105 1.65 4.105 1.03 4.165 1.03 4.165 1.65 5.385 1.65 5.385 1.345 5.505 1.345 5.505 1.405 5.445 1.405 5.445 1.65 6.34 1.65 6.34 1.315 6.4 1.315 6.4 1.65 6.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.8 0.06 6.4 0.06 6.4 0.45 6.34 0.45 6.34 0.06 5.37 0.06 5.37 0.45 5.31 0.45 5.31 0.06 4.145 0.06 4.145 0.29 4.085 0.29 4.085 0.06 3.285 0.06 3.285 0.39 3.165 0.39 3.165 0.33 3.225 0.33 3.225 0.06 1.84 0.06 1.84 0.48 1.9 0.48 1.9 0.54 1.78 0.54 1.78 0.06 1.35 0.06 1.35 0.575 1.29 0.575 1.29 0.06 0.94 0.06 0.94 0.52 0.88 0.52 0.88 0.06 0.575 0.06 0.575 0.2 0.515 0.2 0.515 0.06 0.135 0.06 0.135 0.52 0.075 0.52 0.075 0.06 0 0.06 0 -0.06 6.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.77 1.215 6.605 1.215 6.605 1.34 6.545 1.34 6.545 1.215 6.11 1.215 6.11 0.97 6.05 0.97 6.05 0.91 6.17 0.91 6.17 1.155 6.71 1.155 6.71 0.66 6.605 0.66 6.605 0.355 6.665 0.355 6.665 0.6 6.77 0.6 ;
      POLYGON 6.09 0.475 5.79 0.475 5.79 0.925 5.73 0.925 5.73 1.185 5.985 1.185 5.985 1.34 5.925 1.34 5.925 1.245 4.875 1.245 4.875 1.09 4.745 1.09 4.745 1.03 4.875 1.03 4.875 0.38 4.995 0.38 4.995 0.44 4.935 0.44 4.935 1.185 5.67 1.185 5.67 0.865 5.73 0.865 5.73 0.415 6.03 0.415 6.03 0.355 6.09 0.355 ;
      POLYGON 5.285 1.405 4.585 1.405 4.585 1.29 4.265 1.29 4.265 0.93 4.005 0.93 4.005 1.345 3.34 1.345 3.34 1.285 3.945 1.285 3.945 0.87 4.325 0.87 4.325 1.23 4.585 1.23 4.585 0.87 4.715 0.87 4.715 0.22 5.165 0.22 5.165 0.45 5.105 0.45 5.105 0.28 4.775 0.28 4.775 0.93 4.645 0.93 4.645 1.345 5.285 1.345 ;
      POLYGON 4.615 0.77 4.485 0.77 4.485 1.055 4.425 1.055 4.425 0.77 3.925 0.77 3.925 0.71 4.555 0.71 4.555 0.44 4.495 0.44 4.495 0.38 4.615 0.38 ;
      POLYGON 4.455 0.6 4.335 0.6 4.335 0.45 3.925 0.45 3.925 0.385 3.665 0.385 3.665 0.55 3.605 0.55 3.605 0.735 3.325 0.735 3.325 0.965 3.385 0.965 3.385 1.025 3.265 1.025 3.265 0.735 2.785 0.735 2.785 0.675 2.845 0.675 2.845 0.485 2.905 0.485 2.905 0.675 3.545 0.675 3.545 0.49 3.605 0.49 3.605 0.325 3.985 0.325 3.985 0.39 4.395 0.39 4.395 0.54 4.455 0.54 ;
      POLYGON 4.235 0.61 3.825 0.61 3.825 1.185 2.83 1.185 2.83 0.895 2.625 0.895 2.625 0.475 2.685 0.475 2.685 0.835 2.89 0.835 2.89 1.125 3.765 1.125 3.765 0.485 3.825 0.485 3.825 0.55 4.235 0.55 ;
      POLYGON 2.685 1.15 2.625 1.15 2.625 1.055 1.695 1.055 1.695 0.92 1.655 0.92 1.655 0.8 1.715 0.8 1.715 0.86 1.755 0.86 1.755 0.995 2.465 0.995 2.465 0.595 2.42 0.595 2.42 0.475 2.48 0.475 2.48 0.535 2.525 0.535 2.525 0.995 2.685 0.995 ;
      POLYGON 2.51 1.235 2.005 1.235 2.005 1.3 1.885 1.3 1.885 1.22 1.925 1.22 1.925 1.155 2.51 1.155 ;
      POLYGON 2.135 0.735 1.855 0.735 1.855 0.7 1.555 0.7 1.555 1.09 1.495 1.09 1.495 0.76 1.305 0.76 1.305 0.82 1.245 0.82 1.245 0.7 1.495 0.7 1.495 0.54 1.555 0.54 1.555 0.64 1.915 0.64 1.915 0.675 2.135 0.675 ;
      POLYGON 0.705 1.02 0.625 1.02 0.625 0.85 0.44 0.85 0.44 0.77 0.625 0.77 0.625 0.54 0.705 0.54 ;
  END
END SDFFSX2

MACRO SDFFSX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSX4 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.9814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.74 0.92 7.66 0.92 7.66 0.85 7.505 0.85 7.505 0.715 6.975 0.715 6.975 1.03 6.93 1.03 6.93 1.09 6.87 1.09 6.87 0.97 6.915 0.97 6.915 0.655 7.565 0.655 7.565 0.79 7.74 0.79 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.235 0.815 7.405 1.055 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.61 1.15 6.53 1.15 6.53 0.895 6.365 0.895 6.365 0.815 6.61 0.815 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.43 1.075 6.365 1.075 6.365 1.085 5.94 1.085 5.94 1.005 6.285 1.005 6.285 0.995 6.43 0.995 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 25.04629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.435 0.67 4.375 0.67 4.375 0.42 4.08 0.42 4.08 0.355 3.12 0.355 3.12 0.6 3.14 0.6 3.14 0.73 3.12 0.73 3.12 0.875 2.645 0.875 2.645 0.815 3.06 0.815 3.06 0.295 4.14 0.295 4.14 0.36 4.435 0.36 ;
    END
  END SN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.20925 LAYER Metal1 ;
    ANTENNADIFFAREA 4.620125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4554 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.24297325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 71.231884 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.975 1.405 1.915 1.405 1.915 0.73 1.565 0.73 1.565 1.405 1.505 1.405 1.505 0.73 1.46 0.73 1.46 0.6 1.505 0.6 1.505 0.54 1.565 0.54 1.565 0.67 1.915 0.67 1.915 0.54 1.975 0.54 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.20925 LAYER Metal1 ;
    ANTENNADIFFAREA 4.620125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4554 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.24297325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 71.231884 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.745 1.29 0.685 1.29 0.685 0.92 0.335 0.92 0.335 1.29 0.26 1.29 0.26 0.54 0.335 0.54 0.335 0.79 0.34 0.79 0.34 0.86 0.685 0.86 0.685 0.54 0.745 0.54 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.9 0.13 0.9 0.13 1.65 0.48 1.65 0.48 1.02 0.54 1.02 0.54 1.65 0.89 1.65 0.89 1.17 0.95 1.17 0.95 1.65 1.3 1.65 1.3 1.015 1.36 1.015 1.36 1.65 1.71 1.65 1.71 1.015 1.77 1.015 1.77 1.65 2.12 1.65 2.12 1.095 2.18 1.095 2.18 1.65 2.53 1.65 2.53 1.285 2.59 1.285 2.59 1.65 2.995 1.65 2.995 1.315 3.115 1.315 3.115 1.375 3.055 1.375 3.055 1.65 3.995 1.65 3.995 1.41 4.115 1.41 4.115 1.47 4.055 1.47 4.055 1.65 4.7 1.65 4.7 1.54 4.82 1.54 4.82 1.65 5.94 1.65 5.94 1.51 6 1.51 6 1.65 6.47 1.65 6.47 1.315 6.53 1.315 6.53 1.65 7.375 1.65 7.375 1.315 7.435 1.315 7.435 1.65 8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 0.06 7.45 0.06 7.45 0.555 7.39 0.555 7.39 0.06 6.57 0.06 6.57 0.475 6.51 0.475 6.51 0.06 6.12 0.06 6.12 0.17 6 0.17 6 0.06 4.89 0.06 4.89 0.5 4.83 0.5 4.83 0.06 4.36 0.06 4.36 0.17 4.24 0.17 4.24 0.06 2.62 0.06 2.62 0.49 2.5 0.49 2.5 0.43 2.56 0.43 2.56 0.06 2.18 0.06 2.18 0.52 2.12 0.52 2.12 0.06 1.77 0.06 1.77 0.52 1.71 0.52 1.71 0.06 1.36 0.06 1.36 0.52 1.3 0.52 1.3 0.06 0.98 0.06 0.98 0.2 0.92 0.2 0.92 0.06 0.54 0.06 0.54 0.52 0.48 0.52 0.48 0.06 0.13 0.06 0.13 0.52 0.07 0.52 0.07 0.06 0 0.06 0 -0.06 8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.9 1.215 7.64 1.215 7.64 1.34 7.58 1.34 7.58 1.215 7.075 1.215 7.075 1.06 7.135 1.06 7.135 1.155 7.84 1.155 7.84 0.55 7.565 0.55 7.565 0.49 7.9 0.49 ;
      POLYGON 7.17 0.55 6.785 0.55 6.785 0.635 6.77 0.635 6.77 1.22 6.975 1.22 6.975 1.34 6.915 1.34 6.915 1.28 6.71 1.28 6.71 0.635 6.35 0.635 6.35 0.39 5.84 0.39 5.84 0.38 5.51 0.38 5.51 0.96 5.48 0.96 5.48 1.02 5.42 1.02 5.42 0.9 5.45 0.9 5.45 0.32 5.9 0.32 5.9 0.33 6.41 0.33 6.41 0.575 6.67 0.575 6.67 0.49 7.17 0.49 ;
      POLYGON 6.355 1.31 5.84 1.31 5.84 1.34 4.215 1.34 4.215 1.31 3.62 1.31 3.62 0.9 3.49 0.9 3.49 0.775 3.55 0.775 3.55 0.84 3.68 0.84 3.68 1.25 4.275 1.25 4.275 1.28 5.78 1.28 5.78 0.64 5.84 0.64 5.84 0.49 6.25 0.49 6.25 0.55 5.9 0.55 5.9 0.7 5.84 0.7 5.84 1.25 6.355 1.25 ;
      POLYGON 5.74 0.54 5.68 0.54 5.68 1.18 5.26 1.18 5.26 1.15 3.985 1.15 3.985 0.8 3.94 0.8 3.94 0.68 4 0.68 4 0.74 4.045 0.74 4.045 1.09 5.26 1.09 5.26 0.865 5.245 0.865 5.245 0.73 5.305 0.73 5.305 0.82 5.32 0.82 5.32 1.12 5.62 1.12 5.62 0.48 5.74 0.48 ;
      POLYGON 5.305 0.63 5.145 0.63 5.145 0.93 5.16 0.93 5.16 0.99 5.04 0.99 5.04 0.82 4.695 0.82 4.695 0.76 5.085 0.76 5.085 0.57 5.245 0.57 5.245 0.405 5.305 0.405 ;
      POLYGON 4.985 0.66 4.595 0.66 4.595 0.93 4.655 0.93 4.655 0.99 4.535 0.99 4.535 0.83 4.205 0.83 4.205 0.93 4.265 0.93 4.265 0.99 4.145 0.99 4.145 0.58 3.92 0.58 3.92 0.515 3.795 0.515 3.795 0.455 3.98 0.455 3.98 0.52 4.205 0.52 4.205 0.77 4.535 0.77 4.535 0.6 4.61 0.6 4.61 0.38 4.67 0.38 4.67 0.6 4.985 0.6 ;
      POLYGON 3.885 1.02 3.825 1.02 3.825 0.96 3.78 0.96 3.78 0.74 3.76 0.74 3.76 0.675 3.3 0.675 3.3 1.035 2.485 1.035 2.485 0.915 2.545 0.915 2.545 0.975 3.24 0.975 3.24 0.615 3.525 0.615 3.525 0.455 3.645 0.455 3.645 0.515 3.585 0.515 3.585 0.615 3.82 0.615 3.82 0.68 3.84 0.68 3.84 0.9 3.885 0.9 ;
      POLYGON 3.52 1.105 3.48 1.105 3.48 1.215 2.895 1.215 2.895 1.28 2.775 1.28 2.775 1.2 2.815 1.2 2.815 1.135 3.4 1.135 3.4 1.025 3.52 1.025 ;
      POLYGON 2.94 0.715 2.385 0.715 2.385 1.405 2.325 1.405 2.325 0.76 2.135 0.76 2.135 0.82 2.075 0.82 2.075 0.7 2.325 0.7 2.325 0.485 2.385 0.485 2.385 0.655 2.88 0.655 2.88 0.595 2.94 0.595 ;
      POLYGON 1.155 1.135 1.095 1.135 1.095 0.79 0.845 0.79 0.845 0.73 1.095 0.73 1.095 0.54 1.155 0.54 ;
  END
END SDFFSX4

MACRO SDFFSXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFSXL 0 0 ;
  SIZE 6.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.197 LAYER Metal1 ;
    ANTENNADIFFAREA 3.288925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2106 LAYER Metal1 ;
      ANTENNAMAXAREACAR 15.18043675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 117.22222225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.65 1.16 0.65 1.16 0.995 1.14 0.995 1.14 1.11 1.06 1.11 1.06 0.915 1.08 0.915 1.08 0.57 1.2 0.57 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1524 LAYER Metal1 ;
    ANTENNADIFFAREA 3.288925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2106 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.968661 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 116.12535625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 0.73 0.52 0.73 0.52 1.22 0.46 1.22 0.46 0.63 0.42 0.63 0.42 0.57 0.54 0.57 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.27777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.97 0.705 5.485 0.705 5.485 1.025 5.32 1.025 5.32 0.965 5.425 0.965 5.425 0.645 5.615 0.645 5.615 0.585 5.675 0.585 5.675 0.645 5.835 0.645 5.835 0.625 5.965 0.625 5.965 0.645 5.97 0.645 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.945 1.025 5.755 1.025 5.755 0.895 5.585 0.895 5.585 0.815 5.865 0.815 5.865 0.805 5.945 0.805 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.165 0.705 5.06 0.705 5.06 0.98 4.98 0.98 4.98 0.585 5.165 0.585 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.88 0.96 4.685 0.96 4.685 0.705 4.635 0.705 4.635 0.625 4.765 0.625 4.765 0.88 4.88 0.88 ;
    END
  END CK
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 20.5555555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.15 0.47 2.71 0.47 2.71 0.35 2.165 0.35 2.165 0.875 1.965 0.875 1.965 0.895 1.835 0.895 1.835 0.875 1.715 0.875 1.715 0.815 2.105 0.815 2.105 0.29 2.77 0.29 2.77 0.41 3.09 0.41 3.09 0.35 3.15 0.35 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 0 1.77 0 1.65 0.105 1.65 0.105 1.1 0.165 1.1 0.165 1.65 0.85 1.65 0.85 0.995 0.91 0.995 0.91 1.65 1.555 1.65 1.555 1.305 1.615 1.305 1.615 1.65 1.95 1.65 1.95 1.335 2.07 1.335 2.07 1.395 2.01 1.395 2.01 1.65 3.125 1.65 3.125 1.54 3.245 1.54 3.245 1.65 3.695 1.65 3.695 1.51 3.755 1.51 3.755 1.65 5.03 1.65 5.03 1.285 5.09 1.285 5.09 1.65 5.83 1.65 5.83 1.285 5.89 1.285 5.89 1.65 6.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 5.91 0.06 5.91 0.485 5.85 0.485 5.85 0.06 4.98 0.06 4.98 0.485 4.92 0.485 4.92 0.06 3.79 0.06 3.79 0.41 3.73 0.41 3.73 0.06 2.99 0.06 2.99 0.17 2.87 0.17 2.87 0.06 1.69 0.06 1.69 0.545 1.63 0.545 1.63 0.06 0.88 0.06 0.88 0.2 0.82 0.2 0.82 0.06 0.1 0.06 0.1 0.545 0.16 0.545 0.16 0.605 0.04 0.605 0.04 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.13 1.185 6.095 1.185 6.095 1.31 6.035 1.31 6.035 1.185 5.585 1.185 5.585 1.03 5.645 1.03 5.645 1.125 6.07 1.125 6.07 0.39 6.13 0.39 ;
      POLYGON 5.6 0.485 5.325 0.485 5.325 0.865 5.22 0.865 5.22 1.125 5.46 1.125 5.46 1.31 5.4 1.31 5.4 1.185 4.475 1.185 4.475 0.465 4.595 0.465 4.595 0.525 4.535 0.525 4.535 1.125 5.16 1.125 5.16 0.805 5.265 0.805 5.265 0.425 5.54 0.425 5.54 0.365 5.6 0.365 ;
      POLYGON 4.915 1.345 4.055 1.345 4.055 1.405 3.995 1.405 3.995 1.345 3.595 1.345 3.595 1.37 2.965 1.37 2.965 1.31 3.535 1.31 3.535 1.285 4.315 1.285 4.315 0.305 4.775 0.305 4.775 0.485 4.715 0.485 4.715 0.365 4.375 0.365 4.375 1.285 4.915 1.285 ;
      POLYGON 4.215 1.08 4.155 1.08 4.155 0.89 3.57 0.89 3.57 0.83 4.155 0.83 4.155 0.44 4.215 0.44 ;
      POLYGON 4.055 0.73 3.995 0.73 3.995 0.57 3.57 0.57 3.57 0.44 3.31 0.44 3.31 0.675 3.01 0.675 3.01 1.05 2.89 1.05 2.89 0.99 2.95 0.99 2.95 0.675 2.645 0.675 2.645 0.735 2.585 0.735 2.585 0.615 2.725 0.615 2.725 0.57 2.845 0.57 2.845 0.615 3.25 0.615 3.25 0.38 3.63 0.38 3.63 0.51 4.055 0.51 ;
      POLYGON 3.895 0.73 3.47 0.73 3.47 1.08 3.435 1.08 3.435 1.21 2.705 1.21 2.705 0.895 2.425 0.895 2.425 0.455 2.59 0.455 2.59 0.515 2.485 0.515 2.485 0.835 2.765 0.835 2.765 1.15 3.375 1.15 3.375 1.02 3.41 1.02 3.41 0.54 3.47 0.54 3.47 0.67 3.895 0.67 ;
      POLYGON 2.56 1.15 2.5 1.15 2.5 1.055 1.555 1.055 1.555 0.805 1.615 0.805 1.615 0.995 2.265 0.995 2.265 0.45 2.325 0.45 2.325 0.995 2.56 0.995 ;
      POLYGON 2.385 1.235 1.85 1.235 1.85 1.3 1.73 1.3 1.73 1.22 1.77 1.22 1.77 1.155 2.385 1.155 ;
      POLYGON 2.005 0.705 1.455 0.705 1.455 1.3 1.29 1.3 1.29 1.24 1.395 1.24 1.395 0.47 0.98 0.47 0.98 0.815 0.86 0.815 0.86 0.755 0.92 0.755 0.92 0.41 1.455 0.41 1.455 0.645 2.005 0.645 ;
      POLYGON 0.715 0.89 0.705 0.89 0.705 1.02 0.645 1.02 0.645 0.83 0.655 0.83 0.655 0.47 0.32 0.47 0.32 0.82 0.26 0.82 0.26 0.41 0.715 0.41 ;
  END
END SDFFSXL

MACRO SDFFTRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFTRX1 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.312725 LAYER Metal1 ;
    ANTENNADIFFAREA 3.4753 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2367 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.9954585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 106.9835235 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1 1.33 0.94 1.33 0.94 0.54 0.86 0.54 0.86 0.41 1 0.41 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.312725 LAYER Metal1 ;
    ANTENNADIFFAREA 3.4753 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2367 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.9954585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 106.9835235 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.325 1.29 0.245 1.29 0.245 0.73 0.06 0.73 0.06 0.6 0.245 0.6 0.245 0.54 0.325 0.54 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.14 0.735 5.865 0.735 5.865 0.6 6.06 0.6 6.06 0.43 6.14 0.43 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.765 0.895 5.62 0.895 5.62 0.46 5.7 0.46 5.7 0.815 5.765 0.815 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.52 0.705 5.365 0.705 5.365 0.875 5.19 0.875 5.19 0.625 5.52 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.145 0.92 3.86 0.92 3.86 0.625 3.94 0.625 3.94 0.785 4.145 0.785 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 1.085 1.1 1.085 1.1 1.005 1.285 1.005 1.285 0.77 1.365 0.77 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 1.77 0 1.77 0 1.65 0.47 1.65 0.47 0.995 0.53 0.995 0.53 1.65 1.145 1.65 1.145 1.21 1.205 1.21 1.205 1.65 1.955 1.65 1.955 1.275 2.075 1.275 2.075 1.335 2.015 1.335 2.015 1.65 2.98 1.65 2.98 1.51 3.04 1.51 3.04 1.65 4.075 1.65 4.075 1.18 4.135 1.18 4.135 1.65 5.435 1.65 5.435 1.355 5.495 1.355 5.495 1.65 6.025 1.65 6.025 0.995 6.085 0.995 6.085 1.65 6.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 0.06 5.465 0.06 5.465 0.36 5.405 0.36 5.405 0.06 4.135 0.06 4.135 0.525 4.075 0.525 4.075 0.06 3.07 0.06 3.07 0.17 2.95 0.17 2.95 0.06 2.075 0.06 2.075 0.17 1.955 0.17 1.955 0.06 1.205 0.06 1.205 0.51 1.145 0.51 1.145 0.06 0.56 0.06 0.56 0.2 0.5 0.2 0.5 0.06 0 0.06 0 -0.06 6.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.3 0.895 5.925 0.895 5.925 1.055 5.82 1.055 5.82 1.115 5.42 1.115 5.42 1.255 4.74 1.255 4.74 0.945 4.87 0.945 4.87 0.55 4.81 0.55 4.81 0.43 4.87 0.43 4.87 0.49 4.93 0.49 4.93 1.005 4.8 1.005 4.8 1.195 5.36 1.195 5.36 1.055 5.76 1.055 5.76 0.995 5.865 0.995 5.865 0.835 6.24 0.835 6.24 0.33 5.935 0.33 5.935 0.27 6.3 0.27 ;
      POLYGON 5.26 0.485 5.09 0.485 5.09 0.975 5.26 0.975 5.26 1.095 5.2 1.095 5.2 1.035 5.03 1.035 5.03 0.425 5.2 0.425 5.2 0.325 4.71 0.325 4.71 0.65 4.77 0.65 4.77 0.71 4.71 0.71 4.71 0.845 4.465 0.845 4.465 0.905 4.405 0.905 4.405 0.785 4.65 0.785 4.65 0.265 5.26 0.265 ;
      POLYGON 4.595 1.205 4.535 1.205 4.535 1.08 3.64 1.08 3.64 1.02 3.7 1.02 3.7 0.665 3.67 0.665 3.67 0.435 3.73 0.435 3.73 0.605 3.76 0.605 3.76 1.02 4.245 1.02 4.245 0.625 4.49 0.625 4.49 0.43 4.55 0.43 4.55 0.685 4.305 0.685 4.305 1.02 4.595 1.02 ;
      POLYGON 3.96 1.24 3.48 1.24 3.48 0.605 3.51 0.605 3.51 0.335 2.625 0.335 2.625 0.715 2.565 0.715 2.565 0.275 3.215 0.275 3.215 0.16 3.335 0.16 3.335 0.275 3.93 0.275 3.93 0.525 3.87 0.525 3.87 0.335 3.57 0.335 3.57 0.665 3.54 0.665 3.54 0.765 3.6 0.765 3.6 0.825 3.54 0.825 3.54 1.18 3.96 1.18 ;
      POLYGON 3.41 0.525 3.38 0.525 3.38 1.045 3.32 1.045 3.32 0.855 2.885 0.855 2.885 0.795 3.32 0.795 3.32 0.525 3.29 0.525 3.29 0.465 3.41 0.465 ;
      POLYGON 3.345 1.27 2.675 1.27 2.675 1.34 2.555 1.34 2.555 1.27 2.185 1.27 2.185 1.175 1.465 1.175 1.465 0.53 1.525 0.53 1.525 1.115 2.185 1.115 2.185 0.665 2.305 0.665 2.305 0.725 2.245 0.725 2.245 1.21 3.345 1.21 ;
      POLYGON 3.175 0.695 2.785 0.695 2.785 1.045 2.725 1.045 2.725 0.435 2.785 0.435 2.785 0.635 3.175 0.635 ;
      POLYGON 2.58 1.045 2.52 1.045 2.52 0.875 2.405 0.875 2.405 0.565 2.28 0.565 2.28 0.335 1.88 0.335 1.88 0.33 1.795 0.33 1.795 0.27 1.915 0.27 1.915 0.275 2.34 0.275 2.34 0.505 2.465 0.505 2.465 0.815 2.58 0.815 ;
      POLYGON 2.085 0.685 1.78 0.685 1.78 0.955 1.84 0.955 1.84 1.015 1.72 1.015 1.72 0.49 1.625 0.49 1.625 0.43 1.365 0.43 1.365 0.67 1.16 0.67 1.16 0.81 1.1 0.81 1.1 0.61 1.305 0.61 1.305 0.37 1.685 0.37 1.685 0.43 1.78 0.43 1.78 0.625 2.085 0.625 ;
      POLYGON 0.76 1.02 0.68 1.02 0.68 0.81 0.425 0.81 0.425 0.73 0.68 0.73 0.68 0.54 0.76 0.54 ;
  END
END SDFFTRX1

MACRO SDFFTRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFTRX2 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.46055 LAYER Metal1 ;
    ANTENNADIFFAREA 3.88975 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.302175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.45213875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 88.95507575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.63 1.28 0.63 1.28 0.79 1.34 0.79 1.34 0.92 1.28 0.92 1.28 1.29 1.22 1.29 1.22 0.57 1.34 0.57 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.46055 LAYER Metal1 ;
    ANTENNADIFFAREA 3.88975 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.302175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.45213875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 88.95507575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 0.73 0.72 0.73 0.72 1.29 0.66 1.29 0.66 0.63 0.62 0.63 0.62 0.57 0.74 0.57 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.345 0.73 6.265 0.73 6.265 0.35 6.26 0.35 6.26 0.22 6.34 0.22 6.34 0.27 6.345 0.27 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.165 1.095 6.035 1.095 6.035 1.005 6.085 1.005 6.085 0.645 6.165 0.645 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.935 0.87 5.765 0.87 5.765 0.895 5.605 0.895 5.605 0.645 5.685 0.645 5.685 0.79 5.935 0.79 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.56 0.91 4.34 0.91 4.34 0.965 4.26 0.965 4.26 0.79 4.48 0.79 4.48 0.685 4.56 0.685 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.6 1.74 1.1 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 1.77 0 1.77 0 1.65 0.455 1.65 0.455 0.9 0.515 0.9 0.515 1.65 0.865 1.65 0.865 0.92 0.925 0.92 0.925 1.65 1.425 1.65 1.425 1.02 1.485 1.02 1.485 1.65 2.31 1.65 2.31 1.25 2.43 1.25 2.43 1.31 2.37 1.31 2.37 1.65 3.375 1.65 3.375 1.51 3.435 1.51 3.435 1.65 4.47 1.65 4.47 1.225 4.53 1.225 4.53 1.65 6 1.65 6 1.51 6.06 1.51 6.06 1.65 6.47 1.65 6.47 1.02 6.53 1.02 6.53 1.65 6.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 0.06 6.03 0.06 6.03 0.545 5.97 0.545 5.97 0.06 4.56 0.06 4.56 0.585 4.5 0.585 4.5 0.06 3.48 0.06 3.48 0.17 3.36 0.17 3.36 0.06 2.43 0.06 2.43 0.505 2.31 0.505 2.31 0.445 2.37 0.445 2.37 0.06 1.575 0.06 1.575 0.17 1.455 0.17 1.455 0.06 0.975 0.06 0.975 0.17 0.855 0.17 0.855 0.06 0.475 0.06 0.475 0.2 0.415 0.2 0.415 0.06 0 0.06 0 -0.06 6.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.505 0.92 6.325 0.92 6.325 1.275 5.1 1.275 5.1 1.155 5.285 1.155 5.285 0.585 5.225 0.585 5.225 0.465 5.285 0.465 5.285 0.525 5.345 0.525 5.345 1.215 6.265 1.215 6.265 0.86 6.445 0.86 6.445 0.45 6.505 0.45 ;
      POLYGON 5.825 0.545 5.505 0.545 5.505 0.995 5.825 0.995 5.825 1.115 5.765 1.115 5.765 1.055 5.445 1.055 5.445 0.485 5.765 0.485 5.765 0.365 5.125 0.365 5.125 0.685 5.185 0.685 5.185 0.745 5.125 0.745 5.125 0.905 4.88 0.905 4.88 0.965 4.82 0.965 4.82 0.845 5.065 0.845 5.065 0.305 5.825 0.305 ;
      POLYGON 4.965 0.745 4.72 0.745 4.72 1.065 4.955 1.065 4.955 1.25 4.895 1.25 4.895 1.125 4.155 1.125 4.155 1.155 4.035 1.155 4.035 1.095 4.095 1.095 4.095 0.5 4.155 0.5 4.155 1.065 4.66 1.065 4.66 0.685 4.905 0.685 4.905 0.49 4.965 0.49 ;
      POLYGON 4.355 0.585 4.295 0.585 4.295 0.4 3.995 0.4 3.995 0.75 3.935 0.75 3.935 1.255 4.355 1.255 4.355 1.315 3.875 1.315 3.875 0.69 3.935 0.69 3.935 0.4 3.025 0.4 3.025 0.79 2.965 0.79 2.965 0.34 4.355 0.34 ;
      POLYGON 3.835 0.59 3.775 0.59 3.775 1.185 3.715 1.185 3.715 0.945 3.285 0.945 3.285 0.885 3.715 0.885 3.715 0.53 3.835 0.53 ;
      POLYGON 3.74 1.41 3.15 1.41 3.15 1.425 3.03 1.425 3.03 1.41 2.645 1.41 2.645 1.15 1.84 1.15 1.84 0.57 1.96 0.57 1.96 0.63 1.9 0.63 1.9 1.09 2.645 1.09 2.645 0.825 2.585 0.825 2.585 0.765 2.705 0.765 2.705 1.35 3.74 1.35 ;
      POLYGON 3.57 0.785 3.185 0.785 3.185 1.185 3.125 1.185 3.125 0.53 3.245 0.53 3.245 0.59 3.185 0.59 3.185 0.725 3.57 0.725 ;
      POLYGON 2.98 1.185 2.92 1.185 2.92 1.125 2.805 1.125 2.805 0.665 2.325 0.665 2.325 0.79 2.265 0.79 2.265 0.605 2.805 0.605 2.805 0.5 2.865 0.5 2.865 1.065 2.98 1.065 ;
      POLYGON 2.535 0.985 2.195 0.985 2.195 0.99 2.075 0.99 2.075 0.93 2.105 0.93 2.105 0.47 1.5 0.47 1.5 0.82 1.44 0.82 1.44 0.47 1.04 0.47 1.04 0.82 0.98 0.82 0.98 0.47 0.255 0.47 0.255 0.435 0.195 0.435 0.195 0.375 0.315 0.375 0.315 0.41 2.165 0.41 2.165 0.925 2.535 0.925 ;
      POLYGON 0.56 0.79 0.28 0.79 0.28 1.02 0.22 1.02 0.22 0.63 0.15 0.63 0.15 0.57 0.28 0.57 0.28 0.73 0.56 0.73 ;
  END
END SDFFTRX2

MACRO SDFFTRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFTRX4 0 0 ;
  SIZE 7.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.121 LAYER Metal1 ;
    ANTENNADIFFAREA 4.447425 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4554 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.0491875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 70.13834 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.86 0.545 6.34 0.545 6.34 0.9 6.75 0.9 6.75 1.29 6.69 1.29 6.69 0.96 6.34 0.96 6.34 1.29 6.26 1.29 6.26 0.79 6.27 0.79 6.27 0.485 6.86 0.485 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.121 LAYER Metal1 ;
    ANTENNADIFFAREA 4.447425 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4554 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.0491875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 70.13834 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.93 1.29 5.87 1.29 5.87 0.96 5.52 0.96 5.52 1.29 5.46 1.29 5.46 0.79 5.48 0.79 5.48 0.545 5.33 0.545 5.33 0.485 5.92 0.485 5.92 0.545 5.54 0.545 5.54 0.9 5.93 0.9 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.34 1.005 2.26 1.005 2.26 0.87 2.24 0.87 2.24 0.525 2.32 0.525 2.32 0.79 2.34 0.79 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.14 0.96 2.06 0.96 2.06 0.87 1.995 0.87 1.995 0.525 2.075 0.525 2.075 0.79 2.14 0.79 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.165 0.91 0.87 0.91 0.87 0.815 0.945 0.815 0.945 0.625 1.165 0.625 ;
    END
  END SE
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.77 1.07 0.69 1.07 0.69 0.745 0.635 0.745 0.635 0.625 0.77 0.625 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.375 0.87 0.14 0.87 0.14 0.92 0.06 0.92 0.06 0.79 0.295 0.79 0.295 0.655 0.375 0.655 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.6 1.77 0 1.77 0 1.65 0.315 1.65 0.315 1.02 0.375 1.02 0.375 1.65 0.785 1.65 0.785 1.33 0.845 1.33 0.845 1.65 2.06 1.65 2.06 1.265 2.12 1.265 2.12 1.65 2.76 1.65 2.76 1.285 2.82 1.285 2.82 1.65 3.745 1.65 3.745 1.075 3.805 1.075 3.805 1.65 4.815 1.65 4.815 1.03 4.875 1.03 4.875 1.65 5.255 1.65 5.255 0.97 5.315 0.97 5.315 1.65 5.665 1.65 5.665 1.06 5.725 1.06 5.725 1.65 6.075 1.65 6.075 0.9 6.135 0.9 6.135 1.65 6.485 1.65 6.485 1.06 6.545 1.06 6.545 1.65 6.92 1.65 6.92 1.02 6.98 1.02 6.98 1.65 7.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.6 0.06 7.18 0.06 7.18 0.435 7.12 0.435 7.12 0.06 6.625 0.06 6.625 0.17 6.505 0.17 6.505 0.06 6.155 0.06 6.155 0.17 6.035 0.17 6.035 0.06 5.685 0.06 5.685 0.17 5.565 0.17 5.565 0.06 5.215 0.06 5.215 0.17 5.095 0.17 5.095 0.06 4.745 0.06 4.745 0.55 4.685 0.55 4.685 0.06 3.82 0.06 3.82 0.17 3.7 0.17 3.7 0.06 2.675 0.06 2.675 0.635 2.615 0.635 2.615 0.06 2.12 0.06 2.12 0.425 2.06 0.425 2.06 0.06 0.815 0.06 0.815 0.525 0.755 0.525 0.755 0.06 0 0.06 0 -0.06 7.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.385 0.595 7.29 0.595 7.29 0.92 7.185 0.92 7.185 1.29 7.125 1.29 7.125 0.92 6.85 0.92 6.85 0.77 6.97 0.77 6.97 0.86 7.23 0.86 7.23 0.535 7.325 0.535 7.325 0.455 7.385 0.455 ;
      POLYGON 7.13 0.76 7.07 0.76 7.07 0.67 6.96 0.67 6.96 0.385 4.95 0.385 4.95 0.485 5.205 0.485 5.205 0.76 5.36 0.76 5.36 0.87 5.08 0.87 5.08 1.29 5.02 1.29 5.02 0.87 4.845 0.87 4.845 0.93 4.785 0.93 4.785 0.81 5.145 0.81 5.145 0.545 4.89 0.545 4.89 0.325 7.02 0.325 7.02 0.61 7.13 0.61 ;
      POLYGON 5.045 0.71 4.685 0.71 4.685 1.09 4.36 1.09 4.36 1.03 4.625 1.03 4.625 0.71 4.36 0.71 4.36 0.455 4.42 0.455 4.42 0.65 5.045 0.65 ;
      POLYGON 4.525 0.93 4.465 0.93 4.465 0.87 4.2 0.87 4.2 0.355 3.305 0.355 3.305 0.84 3.335 0.84 3.335 0.9 3.215 0.9 3.215 0.84 3.245 0.84 3.245 0.355 2.985 0.355 2.985 0.475 2.945 0.475 2.945 0.575 2.955 0.575 2.955 1.02 2.895 1.02 2.895 0.635 2.885 0.635 2.885 0.415 2.925 0.415 2.925 0.295 3.48 0.295 3.48 0.215 3.6 0.215 3.6 0.295 4.26 0.295 4.26 0.81 4.525 0.81 ;
      POLYGON 4.1 1.1 4.04 1.1 4.04 0.875 3.65 0.875 3.65 0.815 4.04 0.815 4.04 0.455 4.1 0.455 ;
      POLYGON 3.94 0.715 3.495 0.715 3.495 1.1 3.435 1.1 3.435 0.545 3.405 0.545 3.405 0.485 3.525 0.485 3.525 0.545 3.495 0.545 3.495 0.655 3.94 0.655 ;
      POLYGON 3.24 1.18 2.66 1.18 2.66 1.42 2.22 1.42 2.22 1.165 1.705 1.165 1.705 1.29 1.645 1.29 1.645 1.165 1.615 1.165 1.615 0.36 1.735 0.36 1.735 0.42 1.675 0.42 1.675 1.105 2.28 1.105 2.28 1.36 2.6 1.36 2.6 1.12 3.055 1.12 3.055 0.7 3.085 0.7 3.085 0.455 3.145 0.455 3.145 0.76 3.115 0.76 3.115 1.06 3.24 1.06 ;
      POLYGON 2.795 0.795 2.5 0.795 2.5 1.26 2.38 1.26 2.38 1.2 2.44 1.2 2.44 0.425 2.315 0.425 2.315 0.305 2.375 0.305 2.375 0.365 2.5 0.365 2.5 0.735 2.795 0.735 ;
      POLYGON 1.895 1.005 1.775 1.005 1.775 0.945 1.835 0.945 1.835 0.225 1.08 0.225 1.08 0.465 1.325 0.465 1.325 1.07 0.99 1.07 0.99 1.01 1.265 1.01 1.265 0.525 1.02 0.525 1.02 0.165 1.895 0.165 ;
      POLYGON 1.5 1.29 1.44 1.29 1.44 1.23 0.52 1.23 0.52 0.985 0.475 0.985 0.475 0.52 0.415 0.52 0.415 0.46 0.535 0.46 0.535 0.925 0.58 0.925 0.58 1.17 1.44 1.17 1.44 0.33 1.5 0.33 ;
  END
END SDFFTRX4

MACRO SDFFTRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFTRXL 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.31455 LAYER Metal1 ;
    ANTENNADIFFAREA 3.310925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2106 LAYER Metal1 ;
      ANTENNAMAXAREACAR 15.738604 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 119.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.02 0.57 0.94 0.57 0.94 1.21 0.86 1.21 0.86 0.45 1.02 0.45 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.31455 LAYER Metal1 ;
    ANTENNADIFFAREA 3.310925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2106 LAYER Metal1 ;
      ANTENNAMAXAREACAR 15.738604 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 119.23076925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.305 1.02 0.225 1.02 0.225 0.73 0.06 0.73 0.06 0.6 0.225 0.6 0.225 0.54 0.305 0.54 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.21 0.805 5.865 0.805 5.865 0.725 6.035 0.725 6.035 0.57 6.21 0.57 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.765 0.705 5.545 0.705 5.545 0.905 5.465 0.905 5.465 0.625 5.765 0.625 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.235 0.625 5.365 1.075 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.19 0.91 4.14 0.91 4.14 0.965 4.06 0.965 4.06 0.79 4.11 0.79 4.11 0.515 4.19 0.515 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.37 0.915 1.365 0.915 1.365 1.085 1.04 1.085 1.04 1.005 1.25 1.005 1.25 0.835 1.37 0.835 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 1.77 0 1.77 0 1.65 0.475 1.65 0.475 0.995 0.535 0.995 0.535 1.65 1.17 1.65 1.17 1.185 1.23 1.185 1.23 1.65 2.01 1.65 2.01 1.31 2.13 1.31 2.13 1.37 2.07 1.37 2.07 1.65 3.035 1.65 3.035 1.51 3.095 1.51 3.095 1.65 4.1 1.65 4.1 1.225 4.16 1.225 4.16 1.65 5.31 1.65 5.31 1.35 5.37 1.35 5.37 1.65 5.85 1.65 5.85 1.065 5.91 1.065 5.91 1.65 6.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 0.06 5.455 0.06 5.455 0.5 5.395 0.5 5.395 0.06 4.19 0.06 4.19 0.415 4.13 0.415 4.13 0.06 3.155 0.06 3.155 0.17 3.035 0.17 3.035 0.06 2.13 0.06 2.13 0.17 2.01 0.17 2.01 0.06 1.19 0.06 1.19 0.2 1.13 0.2 1.13 0.06 0.565 0.06 0.565 0.2 0.505 0.2 0.505 0.06 0 0.06 0 -0.06 6.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.37 0.965 5.705 0.965 5.705 1.25 4.73 1.25 4.73 1.005 4.915 1.005 4.915 0.525 4.855 0.525 4.855 0.32 4.915 0.32 4.915 0.465 4.975 0.465 4.975 1.065 4.79 1.065 4.79 1.19 5.645 1.19 5.645 0.905 6.31 0.905 6.31 0.47 5.82 0.47 5.82 0.41 6.37 0.41 ;
      POLYGON 5.25 0.5 5.135 0.5 5.135 1.09 5.075 1.09 5.075 0.44 5.19 0.44 5.19 0.22 4.755 0.22 4.755 0.625 4.815 0.625 4.815 0.685 4.755 0.685 4.755 0.905 4.51 0.905 4.51 0.965 4.45 0.965 4.45 0.845 4.695 0.845 4.695 0.16 5.25 0.16 ;
      POLYGON 4.595 0.745 4.35 0.745 4.35 1.065 4.585 1.065 4.585 1.25 4.525 1.25 4.525 1.125 3.695 1.125 3.695 1.005 3.725 1.005 3.725 0.455 3.785 0.455 3.785 1.065 4.29 1.065 4.29 0.685 4.535 0.685 4.535 0.32 4.595 0.32 ;
      POLYGON 3.985 0.415 3.925 0.415 3.925 0.355 3.625 0.355 3.625 0.685 3.595 0.685 3.595 1.225 3.985 1.225 3.985 1.285 3.535 1.285 3.535 0.625 3.565 0.625 3.565 0.355 2.68 0.355 2.68 0.745 2.62 0.745 2.62 0.295 3.27 0.295 3.27 0.18 3.39 0.18 3.39 0.295 3.985 0.295 ;
      POLYGON 3.465 0.525 3.435 0.525 3.435 1.065 3.375 1.065 3.375 0.875 2.94 0.875 2.94 0.815 3.345 0.815 3.345 0.465 3.465 0.465 ;
      POLYGON 3.4 1.29 3.195 1.29 3.195 1.25 2.73 1.25 2.73 1.38 2.61 1.38 2.61 1.25 2.23 1.25 2.23 1.21 1.465 1.21 1.465 1.09 1.47 1.09 1.47 0.505 1.59 0.505 1.59 0.565 1.53 0.565 1.53 1.15 2.24 1.15 2.24 0.685 2.36 0.685 2.36 0.745 2.3 0.745 2.3 1.19 3.255 1.19 3.255 1.23 3.4 1.23 ;
      POLYGON 3.23 0.715 2.84 0.715 2.84 1.065 2.78 1.065 2.78 0.455 2.84 0.455 2.84 0.655 3.23 0.655 ;
      POLYGON 2.635 1.065 2.575 1.065 2.575 1.005 2.46 1.005 2.46 0.49 1.935 0.49 1.935 0.35 1.85 0.35 1.85 0.29 1.995 0.29 1.995 0.43 2.52 0.43 2.52 0.945 2.635 0.945 ;
      POLYGON 2.14 0.705 1.835 0.705 1.835 0.975 1.895 0.975 1.895 1.035 1.775 1.035 1.775 0.51 1.69 0.51 1.69 0.405 1.185 0.405 1.185 0.735 1.065 0.735 1.065 0.675 1.125 0.675 1.125 0.345 1.75 0.345 1.75 0.45 1.835 0.45 1.835 0.645 2.14 0.645 ;
      POLYGON 0.74 1.02 0.66 1.02 0.66 0.81 0.405 0.81 0.405 0.73 0.66 0.73 0.66 0.54 0.74 0.54 ;
  END
END SDFFTRXL

MACRO SDFFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFX1 0 0 ;
  SIZE 5.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.72865 LAYER Metal1 ;
    ANTENNADIFFAREA 3.0054 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2367 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.5278835 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 88.16856775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 0.73 0.92 0.73 0.92 1.315 0.86 1.315 0.86 0.54 0.92 0.54 0.92 0.6 0.94 0.6 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.77775 LAYER Metal1 ;
    ANTENNADIFFAREA 3.0054 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2367 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.735319 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 89.252218 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.28 1.29 0.2 1.29 0.2 0.73 0.06 0.73 0.06 0.6 0.2 0.6 0.2 0.54 0.28 0.54 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.388889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.165 0.705 4.93 0.705 4.93 0.7 4.44 0.7 4.44 0.965 4.32 0.965 4.32 0.905 4.38 0.905 4.38 0.64 4.93 0.64 4.93 0.585 4.99 0.585 4.99 0.625 5.165 0.625 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.21 0.935 4.76 0.935 4.76 0.855 4.835 0.855 4.835 0.805 5.21 0.805 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.06 0.965 3.98 0.965 3.98 0.73 3.86 0.73 3.86 0.585 3.94 0.585 3.94 0.65 4.06 0.65 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.28 0.96 1.27 0.96 1.27 1.085 1.035 1.085 1.035 1.005 1.19 1.005 1.19 0.88 1.2 0.88 1.2 0.75 1.28 0.75 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 1.77 0 1.77 0 1.65 0.425 1.65 0.425 0.9 0.485 0.9 0.485 1.65 1.065 1.65 1.065 1.195 1.125 1.195 1.125 1.65 1.935 1.65 1.935 1.49 2.055 1.49 2.055 1.55 1.995 1.55 1.995 1.65 2.905 1.65 2.905 1.51 2.965 1.51 2.965 1.65 3.955 1.65 3.955 1.225 4.075 1.225 4.075 1.285 4.015 1.285 4.015 1.65 4.855 1.65 4.855 1.195 4.915 1.195 4.915 1.65 5.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 0.06 4.915 0.06 4.915 0.485 4.855 0.485 4.855 0.06 4.06 0.06 4.06 0.485 4 0.485 4 0.06 2.995 0.06 2.995 0.17 2.875 0.17 2.875 0.06 2.055 0.06 2.055 0.17 1.935 0.17 1.935 0.06 1.095 0.06 1.095 0.43 1.155 0.43 1.155 0.49 1.035 0.49 1.035 0.06 0.515 0.06 0.515 0.2 0.455 0.2 0.455 0.06 0 0.06 0 -0.06 5.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.37 1.095 5.12 1.095 5.12 1.22 5.06 1.22 5.06 1.095 4.6 1.095 4.6 0.86 4.54 0.86 4.54 0.8 4.66 0.8 4.66 1.035 5.31 1.035 5.31 0.525 5.09 0.525 5.09 0.39 5.15 0.39 5.15 0.465 5.37 0.465 ;
      POLYGON 4.605 0.51 4.28 0.51 4.28 0.805 4.22 0.805 4.22 1.065 4.43 1.065 4.43 1.22 4.37 1.22 4.37 1.125 3.625 1.125 3.625 1.185 3.565 1.185 3.565 1.065 3.595 1.065 3.595 0.52 3.655 0.52 3.655 1.065 4.16 1.065 4.16 0.745 4.22 0.745 4.22 0.45 4.545 0.45 4.545 0.39 4.605 0.39 ;
      POLYGON 3.885 0.455 3.755 0.455 3.755 0.42 3.495 0.42 3.495 0.745 3.465 0.745 3.465 1.285 3.725 1.285 3.725 1.225 3.855 1.225 3.855 1.285 3.785 1.285 3.785 1.345 3.405 1.345 3.405 0.685 3.435 0.685 3.435 0.42 2.605 0.42 2.605 0.8 2.545 0.8 2.545 0.36 3.15 0.36 3.15 0.275 3.27 0.275 3.27 0.36 3.815 0.36 3.815 0.395 3.885 0.395 ;
      POLYGON 3.335 0.585 3.305 0.585 3.305 1.15 3.245 1.15 3.245 0.96 2.865 0.96 2.865 0.9 3.215 0.9 3.215 0.525 3.335 0.525 ;
      POLYGON 3.27 1.375 2.615 1.375 2.615 1.425 2.495 1.425 2.495 1.375 2.225 1.375 2.225 1.28 1.37 1.28 1.37 1.02 1.415 1.02 1.415 0.54 1.475 0.54 1.475 1.08 1.43 1.08 1.43 1.22 2.225 1.22 2.225 0.83 2.165 0.83 2.165 0.77 2.285 0.77 2.285 1.315 3.27 1.315 ;
      POLYGON 3.06 0.8 2.765 0.8 2.765 1.12 2.64 1.12 2.64 1.06 2.705 1.06 2.705 0.55 2.825 0.55 2.825 0.61 2.765 0.61 2.765 0.74 3 0.74 3 0.68 3.06 0.68 ;
      POLYGON 2.445 1.15 2.385 1.15 2.385 0.555 1.86 0.555 1.86 0.415 1.775 0.415 1.775 0.355 1.92 0.355 1.92 0.495 2.445 0.495 ;
      POLYGON 2.065 0.77 1.76 0.77 1.76 1.06 1.82 1.06 1.82 1.12 1.7 1.12 1.7 0.575 1.615 0.575 1.615 0.44 1.315 0.44 1.315 0.65 1.1 0.65 1.1 0.82 1.04 0.82 1.04 0.59 1.255 0.59 1.255 0.38 1.675 0.38 1.675 0.515 1.76 0.515 1.76 0.71 2.065 0.71 ;
      POLYGON 0.72 1.02 0.64 1.02 0.64 0.79 0.38 0.79 0.38 0.71 0.64 0.71 0.64 0.54 0.72 0.54 ;
  END
END SDFFX1

MACRO SDFFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFX2 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.08145 LAYER Metal1 ;
    ANTENNADIFFAREA 3.336525 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.302175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.19756775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 79.2752545 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.99 0.63 4.96 0.63 4.96 1.355 4.9 1.355 4.9 0.73 4.86 0.73 4.86 0.6 4.87 0.6 4.87 0.57 4.99 0.57 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.02815 LAYER Metal1 ;
    ANTENNADIFFAREA 3.336525 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.302175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.02117975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 78.3569125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.54 0.73 4.52 0.73 4.52 1.355 4.46 1.355 4.46 0.63 4.4 0.63 4.4 0.57 4.52 0.57 4.52 0.6 4.54 0.6 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.06 0.46 4.14 0.96 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.92 1.26 0.92 1.26 1.21 1.18 1.21 1.18 0.84 1.26 0.84 1.26 0.79 1.34 0.79 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 1.3 0.66 1.3 0.66 1.075 0.44 1.075 0.44 0.995 0.74 0.995 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.787037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 0.895 0.34 0.895 0.34 0.935 0.26 0.935 0.26 0.895 0.235 0.895 0.235 0.815 0.74 0.815 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 0 1.77 0 1.65 0.405 1.65 0.405 1.22 0.465 1.22 0.465 1.65 1.245 1.65 1.245 1.49 1.365 1.49 1.365 1.55 1.305 1.55 1.305 1.65 2.37 1.65 2.37 1.54 2.49 1.54 2.49 1.65 3.325 1.65 3.325 1.49 3.445 1.49 3.445 1.55 3.385 1.55 3.385 1.65 4.255 1.65 4.255 0.965 4.315 0.965 4.315 1.65 4.695 1.65 4.695 0.965 4.755 0.965 4.755 1.65 5.105 1.65 5.105 1.06 5.165 1.06 5.165 1.65 5.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5.195 0.06 5.195 0.2 5.135 0.2 5.135 0.06 4.755 0.06 4.755 0.17 4.635 0.17 4.635 0.06 4.285 0.06 4.285 0.17 4.165 0.17 4.165 0.06 3.355 0.06 3.355 0.52 3.415 0.52 3.415 0.58 3.295 0.58 3.295 0.06 2.485 0.06 2.485 0.17 2.365 0.17 2.365 0.06 1.305 0.06 1.305 0.585 1.245 0.585 1.245 0.06 0.435 0.06 0.435 0.495 0.495 0.495 0.495 0.555 0.375 0.555 0.375 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.425 0.65 5.395 0.65 5.395 1.085 5.315 1.085 5.315 0.915 5.06 0.915 5.06 0.835 5.305 0.835 5.305 0.57 5.425 0.57 ;
      POLYGON 5.415 0.36 4.7 0.36 4.7 0.845 4.64 0.845 4.64 0.36 4.3 0.36 4.3 0.73 4.36 0.73 4.36 0.79 4.24 0.79 4.24 0.36 3.59 0.36 3.59 0.49 3.62 0.49 3.62 1.07 3.68 1.07 3.68 1.13 3.56 1.13 3.56 0.925 3.405 0.925 3.405 0.985 3.345 0.985 3.345 0.865 3.56 0.865 3.56 0.55 3.53 0.55 3.53 0.3 5.415 0.3 ;
      POLYGON 4.065 1.385 2.095 1.385 2.095 1.325 4.005 1.325 4.005 1.12 3.9 1.12 3.9 0.63 3.84 0.63 3.84 0.57 3.96 0.57 3.96 1.06 4.065 1.06 ;
      POLYGON 3.46 0.765 3.245 0.765 3.245 1.145 2.92 1.145 2.92 1.085 3.185 1.085 3.185 0.765 3.135 0.765 3.135 0.605 2.98 0.605 2.98 0.545 3.195 0.545 3.195 0.705 3.46 0.705 ;
      POLYGON 3.085 0.985 3.025 0.985 3.025 0.925 2.82 0.925 2.82 0.81 2.76 0.81 2.76 0.69 2.82 0.69 2.82 0.43 1.925 0.43 1.925 0.835 1.96 0.835 1.96 0.895 1.84 0.895 1.84 0.835 1.865 0.835 1.865 0.43 1.535 0.43 1.535 1.155 1.745 1.155 1.745 1.215 1.475 1.215 1.475 0.37 2.09 0.37 2.09 0.18 2.21 0.18 2.21 0.37 2.88 0.37 2.88 0.865 3.085 0.865 ;
      POLYGON 2.72 0.59 2.66 0.59 2.66 0.91 2.695 0.91 2.695 1.16 2.635 1.16 2.635 0.97 2.275 0.97 2.275 0.91 2.6 0.91 2.6 0.53 2.72 0.53 ;
      POLYGON 2.5 0.765 2.12 0.765 2.12 1.16 2.06 1.16 2.06 0.605 2.025 0.605 2.025 0.545 2.145 0.545 2.145 0.705 2.5 0.705 ;
      POLYGON 1.915 1.375 0.84 1.375 0.84 0.58 0.755 0.58 0.755 0.52 0.9 0.52 0.9 1.315 1.855 1.315 1.855 1.055 1.68 1.055 1.68 0.605 1.645 0.605 1.645 0.545 1.765 0.545 1.765 0.605 1.74 0.605 1.74 0.995 1.915 0.995 ;
      POLYGON 1.06 1.03 1 1.03 1 0.24 0.655 0.24 0.655 0.715 0.135 0.715 0.135 1.035 0.26 1.035 0.26 1.245 0.2 1.245 0.2 1.095 0.075 1.095 0.075 0.655 0.2 0.655 0.2 0.49 0.26 0.49 0.26 0.655 0.595 0.655 0.595 0.18 1.06 0.18 ;
  END
END SDFFX2

MACRO SDFFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFX4 0 0 ;
  SIZE 7 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7802 LAYER Metal1 ;
    ANTENNADIFFAREA 4.307975 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4554 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.3008345 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 64.2028985 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.26 0.55 5.74 0.55 5.74 0.9 6.15 0.9 6.15 1.29 6.09 1.29 6.09 0.96 5.74 0.96 5.74 1.29 5.66 1.29 5.66 0.79 5.67 0.79 5.67 0.49 6.26 0.49 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7802 LAYER Metal1 ;
    ANTENNADIFFAREA 4.307975 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4554 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.3008345 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 64.2028985 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.33 1.29 5.27 1.29 5.27 0.96 4.92 0.96 4.92 1.29 4.86 1.29 4.86 0.79 4.88 0.79 4.88 0.55 4.73 0.55 4.73 0.49 5.32 0.49 5.32 0.55 4.94 0.55 4.94 0.9 5.33 0.9 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.765 0.895 1.635 0.895 1.635 0.72 1.44 0.72 1.44 0.64 1.765 0.64 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.38 1.34 0.88 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.66 1.11 0.54 1.11 0.54 1.17 0.46 1.17 0.46 0.98 0.58 0.98 0.58 0.79 0.66 0.79 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.35185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.84 0.96 0.76 0.96 0.76 0.69 0.34 0.69 0.34 0.73 0.26 0.73 0.26 0.6 0.395 0.6 0.395 0.57 0.475 0.57 0.475 0.6 0.84 0.6 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7 1.77 0 1.77 0 1.65 0.525 1.65 0.525 1.27 0.585 1.27 0.585 1.65 1.37 1.65 1.37 1.3 1.49 1.3 1.49 1.36 1.43 1.36 1.43 1.65 2.245 1.65 2.245 1.54 2.365 1.54 2.365 1.65 3.06 1.65 3.06 1.075 3.12 1.075 3.12 1.65 4.215 1.65 4.215 1.03 4.275 1.03 4.275 1.65 4.655 1.65 4.655 0.97 4.715 0.97 4.715 1.65 5.065 1.65 5.065 1.06 5.125 1.06 5.125 1.65 5.475 1.65 5.475 0.9 5.535 0.9 5.535 1.65 5.885 1.65 5.885 1.06 5.945 1.06 5.945 1.65 6.32 1.65 6.32 1.025 6.38 1.025 6.38 1.65 7 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7 0.06 6.58 0.06 6.58 0.44 6.52 0.44 6.52 0.06 6.025 0.06 6.025 0.17 5.905 0.17 5.905 0.06 5.555 0.06 5.555 0.17 5.435 0.17 5.435 0.06 5.085 0.06 5.085 0.17 4.965 0.17 4.965 0.06 4.615 0.06 4.615 0.17 4.495 0.17 4.495 0.06 4.145 0.06 4.145 0.55 4.085 0.55 4.085 0.06 3.12 0.06 3.12 0.19 3.18 0.19 3.18 0.25 3.06 0.25 3.06 0.06 1.94 0.06 1.94 0.38 1.88 0.38 1.88 0.06 1.415 0.06 1.415 0.28 1.355 0.28 1.355 0.06 0.56 0.06 0.56 0.2 0.5 0.2 0.5 0.06 0 0.06 0 -0.06 7 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.785 0.6 6.69 0.6 6.69 0.925 6.585 0.925 6.585 1.29 6.525 1.29 6.525 0.925 6.25 0.925 6.25 0.77 6.37 0.77 6.37 0.865 6.63 0.865 6.63 0.54 6.725 0.54 6.725 0.46 6.785 0.46 ;
      POLYGON 6.53 0.765 6.47 0.765 6.47 0.67 6.36 0.67 6.36 0.39 4.35 0.39 4.35 0.49 4.605 0.49 4.605 0.77 4.755 0.77 4.755 0.87 4.48 0.87 4.48 1.29 4.42 1.29 4.42 0.87 4.245 0.87 4.245 0.93 4.185 0.93 4.185 0.81 4.545 0.81 4.545 0.55 4.29 0.55 4.29 0.33 6.42 0.33 6.42 0.61 6.53 0.61 ;
      POLYGON 4.445 0.71 4.085 0.71 4.085 1.09 3.76 1.09 3.76 1.03 4.025 1.03 4.025 0.71 3.76 0.71 3.76 0.455 3.82 0.455 3.82 0.65 4.445 0.65 ;
      POLYGON 3.925 0.93 3.865 0.93 3.865 0.87 3.6 0.87 3.6 0.355 3.34 0.355 3.34 0.41 2.9 0.41 2.9 0.345 2.58 0.345 2.58 0.775 2.64 0.775 2.64 0.835 2.52 0.835 2.52 0.345 2.21 0.345 2.21 0.52 2.26 0.52 2.26 1.095 2.435 1.095 2.435 1.155 2.2 1.155 2.2 0.58 2.15 0.58 2.15 0.285 2.705 0.285 2.705 0.16 2.825 0.16 2.825 0.285 2.96 0.285 2.96 0.35 3.28 0.35 3.28 0.295 3.66 0.295 3.66 0.81 3.925 0.81 ;
      POLYGON 3.5 1.1 3.44 1.1 3.44 0.885 2.965 0.885 2.965 0.825 3.44 0.825 3.44 0.455 3.5 0.455 ;
      POLYGON 3.285 0.715 2.8 0.715 2.8 0.815 2.81 0.815 2.81 1.1 2.75 1.1 2.75 0.875 2.74 0.875 2.74 0.545 2.68 0.545 2.68 0.485 2.8 0.485 2.8 0.655 3.285 0.655 ;
      POLYGON 2.605 1.315 2.145 1.315 2.145 1.425 1.705 1.425 1.705 1.2 1 1.2 1 1.295 0.94 1.295 0.94 0.49 0.805 0.49 0.805 0.43 1 0.43 1 1.14 1.765 1.14 1.765 1.365 2.085 1.365 2.085 1.255 2.545 1.255 2.545 0.995 2.36 0.995 2.36 0.455 2.42 0.455 2.42 0.935 2.605 0.935 ;
      POLYGON 2.1 0.74 1.925 0.74 1.925 1.205 1.985 1.205 1.985 1.265 1.865 1.265 1.865 0.54 1.59 0.54 1.59 0.4 1.65 0.4 1.65 0.48 1.925 0.48 1.925 0.68 2.1 0.68 ;
      POLYGON 1.22 1.04 1.1 1.04 1.1 0.325 0.705 0.325 0.705 0.435 0.32 0.435 0.32 0.495 0.16 0.495 0.16 0.83 0.36 0.83 0.36 1.295 0.3 1.295 0.3 0.89 0.1 0.89 0.1 0.435 0.26 0.435 0.26 0.375 0.645 0.375 0.645 0.265 0.73 0.265 0.73 0.195 0.85 0.195 0.85 0.265 1.16 0.265 1.16 0.98 1.22 0.98 ;
  END
END SDFFX4

MACRO SDFFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SDFFXL 0 0 ;
  SIZE 5.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.946825 LAYER Metal1 ;
    ANTENNADIFFAREA 3.0281 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2106 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.99252125 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 106.011396 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.115 0.62 0.94 0.62 0.94 1.21 0.86 1.21 0.86 0.54 1.035 0.54 1.035 0.5 1.115 0.5 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.946825 LAYER Metal1 ;
    ANTENNADIFFAREA 3.0281 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2106 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.99252125 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 106.011396 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.305 1.02 0.225 1.02 0.225 0.635 0.06 0.635 0.06 0.41 0.305 0.41 ;
    END
  END QN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.9074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.385 0.705 4.86 0.705 4.86 0.895 4.84 0.895 4.84 1.01 4.78 1.01 4.78 0.835 4.8 0.835 4.8 0.585 5.105 0.585 5.105 0.625 5.325 0.625 5.325 0.585 5.385 0.585 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.385 0.96 5.235 0.96 5.235 0.895 4.96 0.895 4.96 0.805 5.385 0.805 ;
    END
  END SI
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.52 0.96 4.44 0.96 4.44 0.92 4.34 0.92 4.34 0.96 4.26 0.96 4.26 0.68 4.34 0.68 4.34 0.785 4.52 0.785 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.415 0.96 1.365 0.96 1.365 1.085 1.04 1.085 1.04 1.005 1.285 1.005 1.285 0.88 1.415 0.88 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 1.77 0 1.77 0 1.65 0.475 1.65 0.475 0.995 0.535 0.995 0.535 1.65 1.26 1.65 1.26 1.185 1.32 1.185 1.32 1.65 2.15 1.65 2.15 1.49 2.27 1.49 2.27 1.55 2.21 1.55 2.21 1.65 3.315 1.65 3.315 1.51 3.375 1.51 3.375 1.65 4.43 1.65 4.43 1.22 4.49 1.22 4.49 1.65 5.24 1.65 5.24 1.22 5.3 1.22 5.3 1.65 5.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 0.06 5.34 0.06 5.34 0.485 5.28 0.485 5.28 0.06 4.54 0.06 4.54 0.485 4.48 0.485 4.48 0.06 3.405 0.06 3.405 0.25 3.285 0.25 3.285 0.19 3.345 0.19 3.345 0.06 2.24 0.06 2.24 0.48 2.3 0.48 2.3 0.54 2.18 0.54 2.18 0.06 1.28 0.06 1.28 0.2 1.22 0.2 1.22 0.06 0.565 0.06 0.565 0.2 0.505 0.2 0.505 0.06 0 0.06 0 -0.06 5.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.545 1.245 5.485 1.245 5.485 1.12 5.025 1.12 5.025 1.055 4.965 1.055 4.965 0.995 5.085 0.995 5.085 1.06 5.485 1.06 5.485 0.39 5.545 0.39 ;
      POLYGON 5.03 0.485 4.7 0.485 4.7 0.735 4.68 0.735 4.68 1.155 4.915 1.155 4.915 1.275 4.855 1.275 4.855 1.215 4.62 1.215 4.62 1.12 4.105 1.12 4.105 1.15 3.985 1.15 3.985 1.09 4.045 1.09 4.045 0.505 4.165 0.505 4.165 0.565 4.105 0.565 4.105 1.06 4.62 1.06 4.62 0.675 4.64 0.675 4.64 0.425 4.97 0.425 4.97 0.365 5.03 0.365 ;
      POLYGON 4.335 0.485 4.275 0.485 4.275 0.405 3.945 0.405 3.945 0.725 3.885 0.725 3.885 0.825 3.945 0.825 3.945 0.885 3.885 0.885 3.885 1.25 4.315 1.25 4.315 1.31 3.825 1.31 3.825 0.665 3.885 0.665 3.885 0.405 3.565 0.405 3.565 0.41 3.125 0.41 3.125 0.37 2.865 0.37 2.865 0.69 2.925 0.69 2.925 0.75 2.805 0.75 2.805 0.31 3.185 0.31 3.185 0.35 3.505 0.35 3.505 0.345 3.55 0.345 3.55 0.295 3.67 0.295 3.67 0.345 4.335 0.345 ;
      POLYGON 3.785 0.565 3.725 0.565 3.725 1.18 3.665 1.18 3.665 0.895 3.185 0.895 3.185 0.835 3.665 0.835 3.665 0.505 3.785 0.505 ;
      POLYGON 3.69 1.405 2.485 1.405 2.485 1.31 1.465 1.31 1.465 1.07 1.515 1.07 1.515 0.55 1.635 0.55 1.635 0.61 1.575 0.61 1.575 1.15 1.525 1.15 1.525 1.25 2.485 1.25 2.485 0.86 2.425 0.86 2.425 0.8 2.545 0.8 2.545 1.345 3.69 1.345 ;
      POLYGON 3.51 0.735 3.085 0.735 3.085 1.18 3.025 1.18 3.025 0.59 2.965 0.59 2.965 0.47 3.025 0.47 3.025 0.53 3.085 0.53 3.085 0.675 3.51 0.675 ;
      POLYGON 2.885 1.15 2.645 1.15 2.645 0.7 2.02 0.7 2.02 0.37 1.96 0.37 1.96 0.31 2.08 0.31 2.08 0.64 2.645 0.64 2.645 0.475 2.705 0.475 2.705 1.09 2.885 1.09 ;
      POLYGON 2.325 0.86 1.975 0.86 1.975 1.09 2.035 1.09 2.035 1.15 1.915 1.15 1.915 0.86 1.86 0.86 1.86 0.53 1.8 0.53 1.8 0.45 1.275 0.45 1.275 0.78 1.155 0.78 1.155 0.72 1.215 0.72 1.215 0.39 1.86 0.39 1.86 0.47 1.92 0.47 1.92 0.8 2.325 0.8 ;
      POLYGON 0.74 1.02 0.66 1.02 0.66 0.85 0.405 0.85 0.405 0.77 0.66 0.77 0.66 0.54 0.74 0.54 ;
  END
END SDFFXL

MACRO SEDFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFHQX1 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7501 LAYER Metal1 ;
    ANTENNADIFFAREA 4.256175 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.341775 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.9724235 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 87.2328285 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.605 0.73 3.545 0.73 3.545 1.29 3.485 1.29 3.485 0.73 3.26 0.73 3.26 0.6 3.34 0.6 3.34 0.67 3.545 0.67 3.545 0.54 3.605 0.54 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.26 0.61 6.34 1.11 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.975 0.99 2.835 0.99 2.835 0.895 2.705 0.895 2.705 0.68 2.825 0.68 2.825 0.815 2.975 0.815 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.82838275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.805 0.94 1.725 0.94 1.725 0.705 1.54 0.705 1.54 0.625 1.805 0.625 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.74 0.97 0.475 0.97 0.475 0.655 0.555 0.655 0.555 0.79 0.74 0.79 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.0957095 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.96 0.695 0.9 0.695 0.9 0.555 0.375 0.555 0.375 0.685 0.365 0.685 0.365 0.705 0.235 0.705 0.235 0.625 0.315 0.625 0.315 0.495 0.96 0.495 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 1.77 0 1.77 0 1.65 0.625 1.65 0.625 1.245 0.685 1.245 0.685 1.65 1.445 1.65 1.445 1.19 1.505 1.19 1.505 1.65 2.865 1.65 2.865 1.25 2.925 1.25 2.925 1.65 3.28 1.65 3.28 0.9 3.34 0.9 3.34 1.65 4.005 1.65 4.005 1.105 4.065 1.105 4.065 1.65 4.975 1.65 4.975 1.54 5.095 1.54 5.095 1.65 6.215 1.65 6.215 1.37 6.335 1.37 6.335 1.65 6.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 0.06 6.2 0.06 6.2 0.35 6.14 0.35 6.14 0.06 5.18 0.06 5.18 0.25 5.24 0.25 5.24 0.31 5.12 0.31 5.12 0.06 4.16 0.06 4.16 0.25 4.22 0.25 4.22 0.31 4.1 0.31 4.1 0.06 3.4 0.06 3.4 0.17 3.28 0.17 3.28 0.06 2.755 0.06 2.755 0.42 2.695 0.42 2.695 0.06 1.525 0.06 1.525 0.305 1.585 0.305 1.585 0.365 1.465 0.365 1.465 0.06 0.685 0.06 0.685 0.395 0.625 0.395 0.625 0.06 0 0.06 0 -0.06 6.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.555 1.335 6.435 1.335 6.435 1.27 6.115 1.27 6.115 1.525 5.25 1.525 5.25 1.44 4.625 1.44 4.625 1.45 4.505 1.45 4.505 1.39 4.565 1.39 4.565 1.38 5.31 1.38 5.31 1.465 6.055 1.465 6.055 1.21 6.065 1.21 6.065 0.45 6.3 0.45 6.3 0.315 6.345 0.315 6.345 0.255 6.405 0.255 6.405 0.375 6.36 0.375 6.36 0.51 6.125 0.51 6.125 1.21 6.495 1.21 6.495 1.275 6.555 1.275 ;
      POLYGON 5.995 0.37 5.955 0.37 5.955 1.365 5.535 1.365 5.535 1.26 4.58 1.26 4.58 0.9 4.425 0.9 4.425 0.96 4.365 0.96 4.365 0.84 4.64 0.84 4.64 0.78 4.7 0.78 4.7 0.9 4.64 0.9 4.64 1.2 5.535 1.2 5.535 0.94 5.45 0.94 5.45 0.88 5.595 0.88 5.595 1.305 5.895 1.305 5.895 0.31 5.935 0.31 5.935 0.25 5.995 0.25 ;
      POLYGON 5.795 1.13 5.695 1.13 5.695 1.01 5.735 1.01 5.735 0.47 3.94 0.47 3.94 0.42 3.56 0.42 3.56 0.44 2.975 0.44 2.975 0.58 2.445 0.58 2.445 1.1 2.385 1.1 2.385 0.44 2.445 0.44 2.445 0.52 2.915 0.52 2.915 0.38 3.5 0.38 3.5 0.36 4 0.36 4 0.41 5.795 0.41 ;
      POLYGON 5.62 0.63 5.35 0.63 5.35 1.04 5.435 1.04 5.435 1.1 5.29 1.1 5.29 1 4.96 1 4.96 0.825 5.02 0.825 5.02 0.94 5.29 0.94 5.29 0.57 5.62 0.57 ;
      POLYGON 5.19 0.84 5.13 0.84 5.13 0.725 4.86 0.725 4.86 1.1 4.74 1.1 4.74 1.04 4.8 1.04 4.8 0.63 4.74 0.63 4.74 0.57 4.86 0.57 4.86 0.665 5.19 0.665 ;
      POLYGON 4.64 0.63 4.54 0.63 4.54 0.74 4.265 0.74 4.265 1.06 4.455 1.06 4.455 1.29 4.395 1.29 4.395 1.12 4.205 1.12 4.205 1.005 3.875 1.005 3.875 0.84 3.935 0.84 3.935 0.945 4.205 0.945 4.205 0.68 4.48 0.68 4.48 0.57 4.64 0.57 ;
      POLYGON 4.105 0.845 4.045 0.845 4.045 0.74 3.775 0.74 3.775 1.32 3.715 1.32 3.715 0.82 3.705 0.82 3.705 0.7 3.72 0.7 3.72 0.52 3.84 0.52 3.84 0.58 3.78 0.58 3.78 0.68 4.105 0.68 ;
      POLYGON 3.135 1.15 2.765 1.15 2.765 1.42 1.605 1.42 1.605 1.09 1.38 1.09 1.38 0.79 1.44 0.79 1.44 1.03 1.665 1.03 1.665 1.36 2.705 1.36 2.705 1.09 3.075 1.09 3.075 0.54 3.135 0.54 ;
      POLYGON 2.605 1.26 1.82 1.26 1.82 1.04 1.905 1.04 1.905 0.505 1.845 0.505 1.845 0.445 1.965 0.445 1.965 1.1 1.88 1.1 1.88 1.2 2.225 1.2 2.225 0.675 2.285 0.675 2.285 1.2 2.545 1.2 2.545 0.81 2.605 0.81 ;
      POLYGON 2.21 0.505 2.125 0.505 2.125 1.1 2.065 1.1 2.065 0.445 2.15 0.445 2.15 0.345 1.745 0.345 1.745 0.525 1.12 0.525 1.12 1.095 1.06 1.095 1.06 0.405 1.12 0.405 1.12 0.465 1.685 0.465 1.685 0.285 2.21 0.285 ;
      POLYGON 1.34 0.69 1.28 0.69 1.28 1.255 0.84 1.255 0.84 1.13 0.27 1.13 0.27 1.19 0.21 1.19 0.21 1.13 0.075 1.13 0.075 0.465 0.155 0.465 0.155 0.405 0.215 0.405 0.215 0.525 0.135 0.525 0.135 1.07 0.84 1.07 0.84 0.845 0.96 0.845 0.96 0.905 0.9 0.905 0.9 1.195 1.22 1.195 1.22 0.63 1.34 0.63 ;
  END
END SEDFFHQX1

MACRO SEDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFHQX2 0 0 ;
  SIZE 6.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7683 LAYER Metal1 ;
    ANTENNADIFFAREA 4.439475 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3771 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.99284 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 78.886237 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.265 1.025 3.06 1.025 3.06 0.495 3.185 0.495 3.185 0.575 3.14 0.575 3.14 0.945 3.265 0.945 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.77 0.96 6.48 0.96 6.48 0.67 6.56 0.67 6.56 0.79 6.77 0.79 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.96 1.185 2.88 1.185 2.88 0.92 2.86 0.92 2.86 0.705 2.96 0.705 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.77227725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.625 0.625 1.775 0.895 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.585 0.74 1.085 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.7557755 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.96 0.655 0.9 0.655 0.9 0.485 0.56 0.485 0.56 0.685 0.365 0.685 0.365 0.705 0.235 0.705 0.235 0.625 0.5 0.625 0.5 0.425 0.96 0.425 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.8 1.77 0 1.77 0 1.65 0.625 1.65 0.625 1.36 0.685 1.36 0.685 1.65 1.495 1.65 1.495 1.155 1.555 1.155 1.555 1.65 2.97 1.65 2.97 1.505 2.91 1.505 2.91 1.445 3.03 1.445 3.03 1.65 3.38 1.65 3.38 1.445 3.5 1.445 3.5 1.505 3.44 1.505 3.44 1.65 4.055 1.65 4.055 0.995 4.115 0.995 4.115 1.65 5.07 1.65 5.07 1.54 5.19 1.54 5.19 1.65 6.32 1.65 6.32 1.22 6.38 1.22 6.38 1.65 6.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.8 0.06 6.295 0.06 6.295 0.41 6.235 0.41 6.235 0.06 5.295 0.06 5.295 0.17 5.175 0.17 5.175 0.06 4.195 0.06 4.195 0.355 4.255 0.355 4.255 0.415 4.135 0.415 4.135 0.06 3.42 0.06 3.42 0.17 3.3 0.17 3.3 0.06 2.8 0.06 2.8 0.445 2.74 0.445 2.74 0.06 1.525 0.06 1.525 0.265 1.585 0.265 1.585 0.325 1.465 0.325 1.465 0.06 0.715 0.06 0.715 0.325 0.595 0.325 0.595 0.06 0 0.06 0 -0.06 6.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.615 1.215 6.48 1.215 6.48 1.12 6.22 1.12 6.22 1.405 4.615 1.405 4.615 1.345 6.16 1.345 6.16 1.06 6.32 1.06 6.32 0.57 6.22 0.57 6.22 0.63 6.16 0.63 6.16 0.51 6.44 0.51 6.44 0.315 6.5 0.315 6.5 0.57 6.38 0.57 6.38 1.06 6.54 1.06 6.54 1.155 6.615 1.155 ;
      POLYGON 6.09 0.43 6.06 0.43 6.06 1.245 5.64 1.245 5.64 1.235 4.675 1.235 4.675 0.895 4.435 0.895 4.435 0.835 4.675 0.835 4.675 0.775 4.84 0.775 4.84 0.835 4.735 0.835 4.735 1.175 5.64 1.175 5.64 0.895 5.58 0.895 5.58 0.835 5.7 0.835 5.7 1.185 6 1.185 6 0.37 6.03 0.37 6.03 0.31 6.09 0.31 ;
      POLYGON 5.86 1.085 5.8 1.085 5.8 0.395 4.415 0.395 4.415 0.575 3.975 0.575 3.975 0.395 2.96 0.395 2.96 0.605 2.49 0.605 2.49 1.055 2.43 1.055 2.43 0.465 2.49 0.465 2.49 0.545 2.9 0.545 2.9 0.335 4.035 0.335 4.035 0.515 4.355 0.515 4.355 0.335 5.86 0.335 ;
      POLYGON 5.685 0.555 5.48 0.555 5.48 1.015 5.54 1.015 5.54 1.075 5.42 1.075 5.42 0.915 5.1 0.915 5.1 0.795 5.16 0.795 5.16 0.855 5.42 0.855 5.42 0.495 5.685 0.495 ;
      POLYGON 5.32 0.755 5.26 0.755 5.26 0.695 5 0.695 5 1.055 4.835 1.055 4.835 0.995 4.94 0.995 4.94 0.555 4.795 0.555 4.795 0.495 5 0.495 5 0.635 5.32 0.635 ;
      POLYGON 4.695 0.555 4.575 0.555 4.575 0.735 4.335 0.735 4.335 0.995 4.565 0.995 4.565 1.245 4.505 1.245 4.505 1.055 4.275 1.055 4.275 0.895 3.885 0.895 3.885 0.835 4.275 0.835 4.275 0.675 4.515 0.675 4.515 0.495 4.695 0.495 ;
      POLYGON 4.175 0.735 3.785 0.735 3.785 0.995 3.91 0.995 3.91 1.115 3.85 1.115 3.85 1.055 3.725 1.055 3.725 0.795 3.695 0.795 3.695 0.675 3.755 0.675 3.755 0.495 3.875 0.495 3.875 0.675 4.175 0.675 ;
      POLYGON 3.705 1.345 2.81 1.345 2.81 1.375 1.655 1.375 1.655 1.055 1.43 1.055 1.43 0.93 1.49 0.93 1.49 0.995 1.715 0.995 1.715 1.315 2.75 1.315 2.75 1.285 3.535 1.285 3.535 0.495 3.655 0.495 3.655 0.555 3.595 0.555 3.595 1.225 3.705 1.225 ;
      POLYGON 2.65 1.215 1.815 1.215 1.815 0.995 1.875 0.995 1.875 0.465 1.845 0.465 1.845 0.405 1.965 0.405 1.965 0.465 1.935 0.465 1.935 1.055 1.875 1.055 1.875 1.155 2.27 1.155 2.27 0.635 2.33 0.635 2.33 1.155 2.59 1.155 2.59 0.775 2.65 0.775 ;
      POLYGON 2.255 0.465 2.17 0.465 2.17 1.055 2.11 1.055 2.11 0.405 2.195 0.405 2.195 0.305 1.745 0.305 1.745 0.485 1.12 0.485 1.12 1.18 1.06 1.18 1.06 1.24 1 1.24 1 1.12 1.06 1.12 1.06 0.365 1.12 0.365 1.12 0.425 1.685 0.425 1.685 0.245 2.255 0.245 ;
      POLYGON 1.34 0.69 1.28 0.69 1.28 1.4 0.84 1.4 0.84 1.245 0.45 1.245 0.45 1.305 0.39 1.305 0.39 1.245 0.075 1.245 0.075 0.435 0.34 0.435 0.34 0.375 0.4 0.375 0.4 0.495 0.135 0.495 0.135 1.185 0.84 1.185 0.84 0.96 0.96 0.96 0.96 1.02 0.9 1.02 0.9 1.34 1.22 1.34 1.22 0.63 1.34 0.63 ;
  END
END SEDFFHQX2

MACRO SEDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFHQX4 0 0 ;
  SIZE 8.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.349835 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.97 0.745 7.91 0.745 7.91 0.705 7.13 0.705 7.13 0.89 7.01 0.89 7.01 0.83 7.07 0.83 7.07 0.645 7.635 0.645 7.635 0.625 7.97 0.625 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.81 0.885 7.565 0.885 7.565 0.965 7.39 0.965 7.39 0.805 7.81 0.805 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.82838275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.75 0.94 6.415 0.94 6.415 0.695 6.495 0.695 6.495 0.815 6.75 0.815 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.26 0.71 5.34 1.21 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.16 0.965 5.08 0.965 5.08 0.895 4.835 0.895 4.835 0.775 5.08 0.775 5.08 0.71 5.16 0.71 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.606225 LAYER Metal1 ;
    ANTENNADIFFAREA 5.15165 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.458775 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.04027025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 79.07144025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.745 1.35 0.685 1.35 0.685 0.73 0.335 0.73 0.335 1.35 0.26 1.35 0.26 0.54 0.335 0.54 0.335 0.6 0.34 0.6 0.34 0.67 0.685 0.67 0.685 0.54 0.745 0.54 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.2 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.96 0.13 0.96 0.13 1.65 0.48 1.65 0.48 0.96 0.54 0.96 0.54 1.65 0.89 1.65 0.89 1.04 0.95 1.04 0.95 1.65 1.37 1.65 1.37 1.315 1.43 1.315 1.43 1.65 2.67 1.65 2.67 1.32 2.61 1.32 2.61 1.26 2.73 1.26 2.73 1.65 3.955 1.65 3.955 1.31 3.895 1.31 3.895 1.25 4.015 1.25 4.015 1.65 5.26 1.65 5.26 1.51 5.32 1.51 5.32 1.65 6.76 1.65 6.76 1.24 6.82 1.24 6.82 1.65 7.56 1.65 7.56 1.24 7.62 1.24 7.62 1.65 8.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.2 0.06 7.62 0.06 7.62 0.525 7.56 0.525 7.56 0.06 6.75 0.06 6.75 0.435 6.69 0.435 6.69 0.06 5.34 0.06 5.34 0.39 5.4 0.39 5.4 0.45 5.28 0.45 5.28 0.06 4.04 0.06 4.04 0.52 3.98 0.52 3.98 0.06 2.74 0.06 2.74 0.49 2.62 0.49 2.62 0.43 2.68 0.43 2.68 0.06 1.4 0.06 1.4 0.52 1.34 0.52 1.34 0.06 0.95 0.06 0.95 0.52 0.89 0.52 0.89 0.06 0.54 0.06 0.54 0.52 0.48 0.52 0.48 0.06 0.13 0.06 0.13 0.52 0.07 0.52 0.07 0.06 0 0.06 0 -0.06 8.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 8.13 1.125 8.045 1.125 8.045 1.185 7.985 1.185 7.985 1.125 7.23 1.125 7.23 0.81 7.29 0.81 7.29 1.065 8.07 1.065 8.07 0.43 8.13 0.43 ;
      POLYGON 7.31 0.545 6.91 0.545 6.91 1.04 7.13 1.04 7.13 1.36 7.07 1.36 7.07 1.1 5.98 1.1 5.98 1.16 5.92 1.16 5.92 1.04 6.025 1.04 6.025 0.575 5.91 0.575 5.91 0.515 6.085 0.515 6.085 1.04 6.85 1.04 6.85 0.485 7.25 0.485 7.25 0.425 7.31 0.425 ;
      POLYGON 6.75 0.705 6.595 0.705 6.595 0.595 6.53 0.595 6.53 0.34 5.605 0.34 5.605 0.61 5.12 0.61 5.12 0.4 4.245 0.4 4.245 0.5 4.495 0.5 4.495 1.02 4.435 1.02 4.435 0.56 4.185 0.56 4.185 0.34 5.18 0.34 5.18 0.55 5.545 0.55 5.545 0.28 6.59 0.28 6.59 0.535 6.655 0.535 6.655 0.645 6.75 0.645 ;
      POLYGON 6.585 1.32 5.76 1.32 5.76 0.99 5.6 0.99 5.6 0.87 5.66 0.87 5.66 0.88 5.865 0.88 5.865 0.675 5.925 0.675 5.925 0.94 5.82 0.94 5.82 1.26 6.525 1.26 6.525 1.2 6.585 1.2 ;
      POLYGON 6.43 0.52 6.305 0.52 6.305 0.775 6.185 0.775 6.185 0.695 6.225 0.695 6.225 0.44 6.43 0.44 ;
      POLYGON 5.765 0.77 5.5 0.77 5.5 1.09 5.66 1.09 5.66 1.43 5.6 1.43 5.6 1.15 5.5 1.15 5.5 1.37 4.115 1.37 4.115 1.15 3.345 1.15 3.345 1.31 3.285 1.31 3.285 1.085 3.44 1.085 3.44 0.575 3.38 0.575 3.38 0.515 3.5 0.515 3.5 1.09 4.175 1.09 4.175 1.31 5.44 1.31 5.44 0.71 5.705 0.71 5.705 0.5 5.765 0.5 ;
      POLYGON 5.085 1.185 4.275 1.185 4.275 0.99 3.82 0.99 3.82 0.73 3.88 0.73 3.88 0.93 4.335 0.93 4.335 1.125 4.675 1.125 4.675 0.56 4.96 0.56 4.96 0.5 5.02 0.5 5.02 0.62 4.735 0.62 4.735 1.065 5.085 1.065 ;
      POLYGON 3.855 1.47 2.9 1.47 2.9 1.16 2.51 1.16 2.51 1.32 1.7 1.32 1.7 1.215 1.38 1.215 1.38 1 1.195 1 1.195 1.35 1.135 1.35 1.135 1 1.05 1 1.05 0.79 0.845 0.79 0.845 0.73 1.05 0.73 1.05 0.545 1.135 0.545 1.135 0.485 1.195 0.485 1.195 0.605 1.11 0.605 1.11 0.94 1.38 0.94 1.38 0.88 1.44 0.88 1.44 1.155 1.76 1.155 1.76 1.26 2.45 1.26 2.45 1.1 2.96 1.1 2.96 1.41 3.855 1.41 ;
      POLYGON 3.805 0.63 3.72 0.63 3.72 0.99 3.6 0.99 3.6 0.93 3.66 0.93 3.66 0.57 3.745 0.57 3.745 0.47 3.6 0.47 3.6 0.415 3.28 0.415 3.28 0.985 3.22 0.985 3.22 0.415 2.9 0.415 2.9 0.675 2.955 0.675 2.955 0.795 2.84 0.795 2.84 0.65 2.46 0.65 2.46 0.415 2.14 0.415 2.14 0.765 2.08 0.765 2.08 0.415 1.76 0.415 1.76 0.895 1.7 0.895 1.7 0.355 2.52 0.355 2.52 0.59 2.84 0.59 2.84 0.355 3.66 0.355 3.66 0.41 3.805 0.41 ;
      POLYGON 3.12 1.31 3.06 1.31 3.06 0.97 2.45 0.97 2.45 0.91 3.06 0.91 3.06 0.575 3 0.575 3 0.515 3.12 0.515 ;
      POLYGON 2.74 0.81 2.35 0.81 2.35 1.16 2.29 1.16 2.29 0.575 2.24 0.575 2.24 0.515 2.36 0.515 2.36 0.75 2.74 0.75 ;
      POLYGON 1.98 0.575 1.92 0.575 1.92 1.16 1.86 1.16 1.86 1.055 1.54 1.055 1.54 0.78 1.27 0.78 1.27 0.84 1.21 0.84 1.21 0.72 1.6 0.72 1.6 0.995 1.86 0.995 1.86 0.515 1.98 0.515 ;
  END
END SEDFFHQX4

MACRO SEDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFHQX8 0 0 ;
  SIZE 8.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.6138615 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.61 0.765 8.55 0.765 8.55 0.705 8.035 0.705 8.035 0.695 7.82 0.695 7.82 1.01 7.76 1.01 7.76 0.635 8.035 0.635 8.035 0.625 8.165 0.625 8.165 0.645 8.61 0.645 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.45 1.075 8.37 1.075 8.37 0.895 8.14 0.895 8.14 0.805 8.45 0.805 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.82838275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.26 0.62 7.34 1.12 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.305 0.72 6.165 0.72 6.165 0.95 6.035 0.95 6.035 0.815 6.085 0.815 6.085 0.64 6.305 0.64 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.74 1.125 2.66 1.125 2.66 0.92 2.585 0.92 2.585 0.7 2.74 0.7 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.9905 LAYER Metal1 ;
    ANTENNADIFFAREA 6.0288 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.645525 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.73091675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 61.633554 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.37 0.645 1.325 0.645 1.325 0.9 1.37 0.9 1.37 1.345 1.31 1.345 1.31 0.96 1.265 0.96 1.265 0.8 0.96 0.8 0.96 1.345 0.9 1.345 0.9 0.8 0.55 0.8 0.55 1.345 0.49 1.345 0.49 0.705 0.14 0.705 0.14 1.345 0.08 1.345 0.08 0.73 0.06 0.73 0.06 0.6 0.08 0.6 0.08 0.54 0.14 0.54 0.14 0.645 0.49 0.645 0.49 0.54 0.55 0.54 0.55 0.74 0.9 0.74 0.9 0.54 0.96 0.54 0.96 0.74 1.265 0.74 1.265 0.585 1.31 0.585 1.31 0.525 1.37 0.525 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.8 1.77 0 1.77 0 1.65 0.285 1.65 0.285 0.9 0.345 0.9 0.345 1.65 0.695 1.65 0.695 0.9 0.755 0.9 0.755 1.65 1.105 1.65 1.105 0.9 1.165 0.9 1.165 1.65 1.515 1.65 1.515 0.955 1.575 0.955 1.575 1.65 1.925 1.65 1.925 1.09 1.985 1.09 1.985 1.65 2.7 1.65 2.7 1.51 2.76 1.51 2.76 1.65 4.16 1.65 4.16 1.25 4.28 1.25 4.28 1.31 4.22 1.31 4.22 1.65 5.64 1.65 5.64 1.51 5.7 1.51 5.7 1.65 6.05 1.65 6.05 1.21 6.17 1.21 6.17 1.27 6.11 1.27 6.11 1.65 7.41 1.65 7.41 1.54 7.53 1.54 7.53 1.65 8.195 1.65 8.195 1.35 8.255 1.35 8.255 1.65 8.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.8 0.06 8.365 0.06 8.365 0.475 8.305 0.475 8.305 0.06 7.44 0.06 7.44 0.27 7.5 0.27 7.5 0.33 7.38 0.33 7.38 0.06 6.255 0.06 6.255 0.38 6.195 0.38 6.195 0.06 5.615 0.06 5.615 0.28 5.555 0.28 5.555 0.06 4.19 0.06 4.19 0.32 4.25 0.32 4.25 0.38 4.13 0.38 4.13 0.06 3.015 0.06 3.015 0.28 2.895 0.28 2.895 0.22 2.955 0.22 2.955 0.06 1.985 0.06 1.985 0.52 1.925 0.52 1.925 0.06 1.575 0.06 1.575 0.52 1.515 0.52 1.515 0.06 1.165 0.06 1.165 0.485 1.105 0.485 1.105 0.06 0.755 0.06 0.755 0.485 0.695 0.485 0.695 0.06 0.345 0.06 0.345 0.485 0.285 0.485 0.285 0.06 0 0.06 0 -0.06 8.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 8.77 1.235 8.49 1.235 8.49 1.295 8.43 1.295 8.43 1.235 7.98 1.235 7.98 1.01 7.92 1.01 7.92 0.95 8.04 0.95 8.04 1.175 8.71 1.175 8.71 0.5 8.625 0.5 8.625 0.38 8.685 0.38 8.685 0.44 8.77 0.44 ;
      POLYGON 8.055 0.5 7.66 0.5 7.66 1.11 7.88 1.11 7.88 1.47 7.82 1.47 7.82 1.17 7.6 1.17 7.6 0.52 7.09 0.52 7.09 1 6.81 1 6.81 0.94 7.03 0.94 7.03 0.52 6.935 0.52 6.935 0.4 6.995 0.4 6.995 0.46 7.6 0.46 7.6 0.44 7.995 0.44 7.995 0.38 8.055 0.38 ;
      POLYGON 7.5 1.44 6.27 1.44 6.27 1.11 5.935 1.11 5.935 1.3 5.875 1.3 5.875 0.4 5.935 0.4 5.935 1.05 6.33 1.05 6.33 1.38 7.44 1.38 7.44 0.91 7.5 0.91 ;
      POLYGON 7.295 1.28 6.65 1.28 6.65 0.79 6.565 0.79 6.565 0.73 6.775 0.73 6.775 0.24 7.265 0.24 7.265 0.36 7.205 0.36 7.205 0.3 6.835 0.3 6.835 0.62 6.93 0.62 6.93 0.74 6.835 0.74 6.835 0.79 6.71 0.79 6.71 1.22 7.295 1.22 ;
      POLYGON 6.675 0.54 6.465 0.54 6.465 0.89 6.49 0.89 6.49 0.94 6.55 0.94 6.55 1 6.43 1 6.43 0.95 6.405 0.95 6.405 0.54 6.035 0.54 6.035 0.3 5.775 0.3 5.775 0.44 5.395 0.44 5.395 0.32 4.86 0.32 4.86 0.58 5.08 0.58 5.08 1.02 5.02 1.02 5.02 0.64 4.8 0.64 4.8 0.26 5.455 0.26 5.455 0.38 5.715 0.38 5.715 0.24 6.095 0.24 6.095 0.48 6.615 0.48 6.615 0.4 6.675 0.4 ;
      POLYGON 5.775 1.34 4.38 1.34 4.38 1.15 4.06 1.15 4.06 1.34 2.86 1.34 2.86 1.285 2.19 1.285 2.19 1.345 2.13 1.345 2.13 0.99 1.78 0.99 1.78 1.345 1.72 1.345 1.72 0.8 1.425 0.8 1.425 0.74 1.72 0.74 1.72 0.54 1.78 0.54 1.78 0.93 2.245 0.93 2.245 0.54 2.305 0.54 2.305 0.99 2.19 0.99 2.19 1.225 2.84 1.225 2.84 0.74 2.9 0.74 2.9 1.235 2.92 1.235 2.92 1.28 4 1.28 4 1.09 4.44 1.09 4.44 1.28 5.715 1.28 5.715 0.74 5.775 0.74 ;
      POLYGON 5.295 1.18 4.54 1.18 4.54 0.99 3.9 0.99 3.9 1.18 3.02 1.18 3.02 0.74 3.08 0.74 3.08 1.12 3.52 1.12 3.52 0.61 3.58 0.61 3.58 1.12 3.84 1.12 3.84 0.93 4.48 0.93 4.48 0.7 4.42 0.7 4.42 0.64 4.54 0.64 4.54 0.93 4.6 0.93 4.6 1.12 4.86 1.12 4.86 0.74 4.92 0.74 4.92 1.12 5.235 1.12 5.235 0.48 5.175 0.48 5.175 0.42 5.295 0.42 ;
      POLYGON 4.76 1.02 4.7 1.02 4.7 0.83 4.64 0.83 4.64 0.54 4.155 0.54 4.155 0.655 4.095 0.655 4.095 0.48 4.495 0.48 4.495 0.375 4.555 0.375 4.555 0.48 4.7 0.48 4.7 0.77 4.76 0.77 ;
      POLYGON 4.325 0.815 3.74 0.815 3.74 1.02 3.68 1.02 3.68 0.375 3.74 0.375 3.74 0.755 4.325 0.755 ;
      POLYGON 3.42 1.02 3.36 1.02 3.36 0.44 2.735 0.44 2.735 0.28 2.145 0.28 2.145 0.83 2.085 0.83 2.085 0.22 2.795 0.22 2.795 0.38 3.36 0.38 3.36 0.32 3.42 0.32 ;
      POLYGON 3.26 0.66 3.2 0.66 3.2 0.6 2.485 0.6 2.485 1.02 2.425 1.02 2.425 0.38 2.635 0.38 2.635 0.44 2.485 0.44 2.485 0.54 3.26 0.54 ;
  END
END SEDFFHQX8

MACRO SEDFFTRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFTRX1 0 0 ;
  SIZE 8.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.580075 LAYER Metal1 ;
    ANTENNADIFFAREA 4.598125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3177 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.416352 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 113.70632675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.54 0.73 5.5 0.73 5.5 1.08 5.315 1.08 5.315 1 5.42 1 5.42 0.54 5.5 0.54 5.5 0.6 5.54 0.6 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.636875 LAYER Metal1 ;
    ANTENNADIFFAREA 4.598125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3177 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.595137 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 114.42870625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.54 0.14 1.29 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.97 1.06 7.94 1.06 7.94 1.17 7.86 1.17 7.86 0.98 7.89 0.98 7.89 0.7 7.97 0.7 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.52777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.54 0.92 7.46 0.92 7.46 0.85 6.985 0.85 6.985 0.77 7.54 0.77 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.11 0.955 5.94 0.955 5.94 1.205 5.86 1.205 5.86 0.875 6.11 0.875 ;
    END
  END RN
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.34 0.92 4.16 0.92 4.16 0.96 4.08 0.96 4.08 0.64 4.34 0.64 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.37962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.66 0.82 4.6 0.82 4.6 0.54 3.98 0.54 3.98 0.82 3.92 0.82 3.92 0.705 3.835 0.705 3.835 0.625 3.92 0.625 3.92 0.48 4.66 0.48 ;
    END
  END SE
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.67 3.35 1.12 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.2 1.77 0 1.77 0 1.65 0.285 1.65 0.285 0.9 0.345 0.9 0.345 1.65 1.015 1.65 1.015 1.34 1.135 1.34 1.135 1.4 1.075 1.4 1.075 1.65 2.1 1.65 2.1 1.28 2.04 1.28 2.04 1.22 2.16 1.22 2.16 1.65 3.165 1.65 3.165 1.54 3.285 1.54 3.285 1.65 4.05 1.65 4.05 1.54 4.17 1.54 4.17 1.65 5.08 1.65 5.08 1.34 5.2 1.34 5.2 1.4 5.14 1.4 5.14 1.65 5.965 1.65 5.965 1.54 6.085 1.54 6.085 1.65 7.875 1.65 7.875 1.43 7.935 1.43 7.935 1.65 8.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.2 0.06 7.905 0.06 7.905 0.6 7.845 0.6 7.845 0.06 6.915 0.06 6.915 0.29 6.975 0.29 6.975 0.35 6.855 0.35 6.855 0.06 6.685 0.06 6.685 0.29 6.745 0.29 6.745 0.35 6.625 0.35 6.625 0.06 6.2 0.06 6.2 0.455 6.08 0.455 6.08 0.395 6.14 0.395 6.14 0.06 5.16 0.06 5.16 0.52 5.1 0.52 5.1 0.06 4.055 0.06 4.055 0.16 4.115 0.16 4.115 0.22 3.995 0.22 3.995 0.06 3.225 0.06 3.225 0.41 3.165 0.41 3.165 0.06 2.16 0.06 2.16 0.25 2.04 0.25 2.04 0.19 2.1 0.19 2.1 0.06 1.125 0.06 1.125 0.635 1.065 0.635 1.065 0.06 0.345 0.06 0.345 0.52 0.285 0.52 0.285 0.06 0 0.06 0 -0.06 8.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 8.13 1.33 7.16 1.33 7.16 1.27 8.07 1.27 8.07 0.505 8.13 0.505 ;
      POLYGON 7.7 1.02 7.64 1.02 7.64 0.67 6.535 0.67 6.535 0.61 7.64 0.61 7.64 0.505 7.7 0.505 ;
      POLYGON 7.31 1.105 7.25 1.105 7.25 1.01 6.9 1.01 6.9 1.105 6.825 1.105 6.825 0.83 6.375 0.83 6.375 0.615 5.92 0.615 5.92 0.32 5.32 0.32 5.32 0.68 5.055 0.68 5.055 0.82 4.995 0.82 4.995 0.62 5.26 0.62 5.26 0.26 5.98 0.26 5.98 0.555 6.315 0.555 6.315 0.39 6.375 0.39 6.375 0.45 7.165 0.45 7.165 0.315 7.285 0.315 7.285 0.375 7.225 0.375 7.225 0.51 6.435 0.51 6.435 0.77 6.885 0.77 6.885 0.95 7.31 0.95 ;
      POLYGON 7.135 1.17 7.06 1.17 7.06 1.295 6.46 1.295 6.46 1.23 6.435 1.23 6.435 1.11 6.495 1.11 6.495 1.175 6.52 1.175 6.52 1.235 7 1.235 7 1.11 7.135 1.11 ;
      POLYGON 6.7 1.135 6.62 1.135 6.62 1.01 6.31 1.01 6.31 1.135 6.23 1.135 6.23 0.93 6.7 0.93 ;
      POLYGON 6.36 1.365 5.3 1.365 5.3 1.24 4.98 1.24 4.98 1.44 2.26 1.44 2.26 1.12 1.94 1.12 1.94 1.375 1.355 1.375 1.355 1.44 1.235 1.44 1.235 1.24 0.565 1.24 0.565 1.245 0.445 1.245 0.445 1.185 0.505 1.185 0.505 1.18 0.84 1.18 0.84 0.54 0.9 0.54 0.9 1.18 1.295 1.18 1.295 1.315 1.88 1.315 1.88 1.06 2.32 1.06 2.32 1.38 4.92 1.38 4.92 1.18 5.155 1.18 5.155 0.84 5.215 0.84 5.215 0.78 5.275 0.78 5.275 0.9 5.215 0.9 5.215 1.18 5.36 1.18 5.36 1.305 6.36 1.305 ;
      POLYGON 6.18 0.775 5.76 0.775 5.76 1.135 5.7 1.135 5.7 0.42 5.82 0.42 5.82 0.48 5.76 0.48 5.76 0.715 6.18 0.715 ;
      POLYGON 4.915 0.255 4.275 0.255 4.275 0.38 3.735 0.38 3.735 1.06 4.44 1.06 4.44 0.78 4.5 0.78 4.5 1.12 3.675 1.12 3.675 0.32 4.215 0.32 4.215 0.195 4.915 0.195 ;
      POLYGON 4.82 0.98 4.66 0.98 4.66 1.28 2.74 1.28 2.74 0.54 2.8 0.54 2.8 1.22 4.6 1.22 4.6 0.92 4.76 0.92 4.76 0.53 4.82 0.53 ;
      POLYGON 3.51 1.02 3.45 1.02 3.45 0.57 3.16 0.57 3.16 0.63 3.1 0.63 3.1 0.51 3.45 0.51 3.45 0.315 3.51 0.315 ;
      POLYGON 3 1.02 2.94 1.02 2.94 0.375 2.64 0.375 2.64 0.95 2.58 0.95 2.58 0.375 2.32 0.375 2.32 0.41 1.385 0.41 1.385 0.86 1.46 0.86 1.46 0.92 1.325 0.92 1.325 0.35 1.625 0.35 1.625 0.34 1.745 0.34 1.745 0.35 2.26 0.35 2.26 0.315 3 0.315 ;
      POLYGON 2.48 1.215 2.42 1.215 2.42 0.8 1.935 0.8 1.935 0.74 2.42 0.74 2.42 0.54 2.48 0.54 ;
      POLYGON 2.265 0.96 1.78 0.96 1.78 1.215 1.72 1.215 1.72 0.54 1.78 0.54 1.78 0.9 2.265 0.9 ;
      POLYGON 1.62 1.215 1.515 1.215 1.515 1.08 1 1.08 1 0.91 1.06 0.91 1.06 1.02 1.56 1.02 1.56 0.63 1.485 0.63 1.485 0.57 1.62 0.57 ;
      POLYGON 0.58 1.02 0.5 1.02 0.5 0.79 0.24 0.79 0.24 0.71 0.5 0.71 0.5 0.54 0.58 0.54 ;
  END
END SEDFFTRX1

MACRO SEDFFTRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFTRX2 0 0 ;
  SIZE 8.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.66055 LAYER Metal1 ;
    ANTENNADIFFAREA 4.90835 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.383175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.16298025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 95.12624775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.19 0.6 5.065 0.6 5.065 1.02 4.985 1.02 4.985 0.73 4.86 0.73 4.86 0.6 4.985 0.6 4.985 0.52 5.19 0.52 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.66055 LAYER Metal1 ;
    ANTENNADIFFAREA 4.90835 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.383175 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.16298025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 95.12624775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.74 0.92 4.685 0.92 4.685 0.99 4.615 0.99 4.615 1.02 4.535 1.02 4.535 0.885 4.6 0.885 4.6 0.52 4.72 0.52 4.72 0.6 4.68 0.6 4.68 0.79 4.74 0.79 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.965 1.065 7.835 1.065 7.835 0.615 7.955 0.615 7.955 0.815 7.965 0.815 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.575 0.895 7.035 0.895 7.035 0.815 7.495 0.815 7.495 0.775 7.575 0.775 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.76 0.815 6.025 1.13 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.26 0.68 4.34 1.18 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.68 0.895 0.19 0.895 0.19 0.805 0.67 0.805 0.67 0.815 0.68 0.815 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 18.37962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.16 0.85 1.1 0.85 1.1 0.36 0.695 0.36 0.695 0.645 0.84 0.645 0.84 0.705 0.235 0.705 0.235 0.625 0.435 0.625 0.435 0.645 0.635 0.645 0.635 0.3 1.16 0.3 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.2 1.77 0 1.77 0 1.65 0.475 1.65 0.475 1.155 0.595 1.155 0.595 1.215 0.535 1.215 0.535 1.65 1.335 1.65 1.335 1.54 1.455 1.54 1.455 1.65 2.26 1.65 2.26 1.51 2.32 1.51 2.32 1.65 3.66 1.65 3.66 1.54 3.78 1.54 3.78 1.65 4.3 1.65 4.3 1.51 4.36 1.51 4.36 1.65 4.74 1.65 4.74 1.46 4.86 1.46 4.86 1.52 4.8 1.52 4.8 1.65 5.24 1.65 5.24 1.51 5.3 1.51 5.3 1.65 6.125 1.65 6.125 1.45 6.065 1.45 6.065 1.39 6.185 1.39 6.185 1.65 7.76 1.65 7.76 1.51 7.82 1.51 7.82 1.65 8.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.2 0.06 7.86 0.06 7.86 0.515 7.8 0.515 7.8 0.06 6.935 0.06 6.935 0.335 6.995 0.335 6.995 0.395 6.875 0.395 6.875 0.06 6.765 0.06 6.765 0.395 6.705 0.395 6.705 0.06 6.17 0.06 6.17 0.17 6.05 0.17 6.05 0.06 5.425 0.06 5.425 0.17 5.305 0.17 5.305 0.06 4.955 0.06 4.955 0.17 4.835 0.17 4.835 0.06 4.485 0.06 4.485 0.17 4.365 0.17 4.365 0.06 3.675 0.06 3.675 0.45 3.735 0.45 3.735 0.51 3.615 0.51 3.615 0.06 2.54 0.06 2.54 0.31 2.42 0.31 2.42 0.25 2.48 0.25 2.48 0.06 1.355 0.06 1.355 0.525 1.295 0.525 1.295 0.06 0.535 0.06 0.535 0.525 0.475 0.525 0.475 0.06 0 0.06 0 -0.06 8.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 8.125 1.235 7.815 1.235 7.815 1.375 7.245 1.375 7.245 1.315 7.755 1.315 7.755 1.175 8.065 1.175 8.065 0.515 8.005 0.515 8.005 0.395 8.065 0.395 8.065 0.455 8.125 0.455 ;
      POLYGON 7.735 1.055 7.655 1.055 7.655 1.14 7.595 1.14 7.595 0.995 7.675 0.995 7.675 0.675 7.595 0.675 7.595 0.435 7.155 0.435 7.155 0.555 6.71 0.555 6.71 0.83 6.65 0.83 6.65 0.495 7.095 0.495 7.095 0.375 7.655 0.375 7.655 0.615 7.735 0.615 ;
      POLYGON 7.395 1.15 7.335 1.15 7.335 1.055 6.985 1.055 6.985 1.15 6.875 1.15 6.875 1.08 6.185 1.08 6.185 1.29 5.965 1.29 5.965 1.515 5.44 1.515 5.44 1.36 4.64 1.36 4.64 1.41 3.56 1.41 3.56 1.47 2.42 1.47 2.42 1.375 1.235 1.375 1.235 1.35 1.175 1.35 1.175 1.29 1.295 1.29 1.295 1.315 2.48 1.315 2.48 1.41 3.5 1.41 3.5 1.35 4.58 1.35 4.58 1.3 5.5 1.3 5.5 1.455 5.905 1.455 5.905 1.23 6.125 1.23 6.125 1.02 6.365 1.02 6.365 0.63 6.285 0.63 6.285 0.57 6.425 0.57 6.425 1.02 6.875 1.02 6.875 0.655 7.255 0.655 7.255 0.535 7.375 0.535 7.375 0.595 7.315 0.595 7.315 0.715 6.935 0.715 6.935 0.995 7.395 0.995 ;
      POLYGON 7.22 1.215 7.145 1.215 7.145 1.31 6.975 1.31 6.975 1.515 6.52 1.515 6.52 1.36 6.58 1.36 6.58 1.455 6.915 1.455 6.915 1.25 7.085 1.25 7.085 1.155 7.22 1.155 ;
      POLYGON 6.815 1.355 6.68 1.355 6.68 1.26 6.405 1.26 6.405 1.355 6.285 1.355 6.285 1.275 6.325 1.275 6.325 1.18 6.76 1.18 6.76 1.275 6.815 1.275 ;
      POLYGON 6.48 0.395 4.5 0.395 4.5 0.77 4.44 0.77 4.44 0.395 3.955 0.395 3.955 0.99 3.5 0.99 3.5 0.93 3.895 0.93 3.895 0.335 5.525 0.335 5.525 0.325 5.645 0.325 5.645 0.335 6.48 0.335 ;
      POLYGON 6.265 0.815 6.125 0.815 6.125 0.715 5.66 0.715 5.66 1.295 5.805 1.295 5.805 1.355 5.6 1.355 5.6 0.655 5.845 0.655 5.845 0.54 5.905 0.54 5.905 0.655 6.185 0.655 6.185 0.755 6.265 0.755 ;
      POLYGON 5.66 0.555 5.5 0.555 5.5 1.02 5.44 1.02 5.44 0.83 5.165 0.83 5.165 0.77 5.44 0.77 5.44 0.495 5.66 0.495 ;
      POLYGON 4.25 0.58 4.125 0.58 4.125 1.15 3.4 1.15 3.4 1.31 2.58 1.31 2.58 1.215 2.2 1.215 2.2 0.9 2.26 0.9 2.26 1.155 2.64 1.155 2.64 1.25 2.96 1.25 2.96 0.93 3.08 0.93 3.08 0.99 3.02 0.99 3.02 1.25 3.34 1.25 3.34 0.77 3.46 0.77 3.46 0.83 3.4 0.83 3.4 1.09 4.065 1.09 4.065 0.52 4.25 0.52 ;
      POLYGON 3.795 0.83 3.735 0.83 3.735 0.67 3.24 0.67 3.24 1.15 3.12 1.15 3.12 1.09 3.18 1.09 3.18 0.54 3.24 0.54 3.24 0.61 3.795 0.61 ;
      POLYGON 3.08 0.82 3.02 0.82 3.02 0.47 2.26 0.47 2.26 0.44 1.94 0.44 1.94 0.95 1.88 0.95 1.88 0.44 1.56 0.44 1.56 0.995 1.62 0.995 1.62 1.055 1.5 1.055 1.5 0.38 2.145 0.38 2.145 0.275 2.265 0.275 2.265 0.38 2.32 0.38 2.32 0.41 3.08 0.41 ;
      POLYGON 2.92 0.63 2.86 0.63 2.86 1.15 2.74 1.15 2.74 1.09 2.8 1.09 2.8 0.99 2.36 0.99 2.36 0.93 2.8 0.93 2.8 0.57 2.92 0.57 ;
      POLYGON 2.635 0.79 2.1 0.79 2.1 1.18 2.04 1.18 2.04 0.57 2.16 0.57 2.16 0.63 2.1 0.63 2.1 0.73 2.635 0.73 ;
      POLYGON 1.875 1.215 1.37 1.215 1.37 1.19 0.94 1.19 0.94 0.52 0.795 0.52 0.795 0.46 1 0.46 1 1.13 1.425 1.13 1.425 1.155 1.72 1.155 1.72 0.54 1.78 0.54 1.78 1.095 1.875 1.095 ;
      POLYGON 0.84 1.055 0.33 1.055 0.33 1.115 0.27 1.115 0.27 1.055 0.03 1.055 0.03 0.465 0.27 0.465 0.27 0.405 0.33 0.405 0.33 0.525 0.09 0.525 0.09 0.995 0.78 0.995 0.78 0.805 0.84 0.805 ;
  END
END SEDFFTRX2

MACRO SEDFFTRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFTRX4 0 0 ;
  SIZE 9.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.352275 LAYER Metal1 ;
    ANTENNADIFFAREA 6.188375 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.5364 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.97814125 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 77.852349 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.425 0.55 5.965 0.55 5.965 1.005 6.17 1.005 6.17 1.025 6.295 1.025 6.295 1.085 6.11 1.085 6.11 1.065 5.965 1.065 5.965 1.085 5.705 1.085 5.705 1.025 5.835 1.025 5.835 1.005 5.905 1.005 5.905 0.55 5.835 0.55 5.835 0.49 6.425 0.49 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.352275 LAYER Metal1 ;
    ANTENNADIFFAREA 6.188375 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.5364 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.97814125 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 77.852349 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.485 0.52 5.12 0.52 5.12 1.005 5.325 1.005 5.325 1.125 5.265 1.125 5.265 1.065 5.165 1.065 5.165 1.085 4.735 1.085 4.735 1.025 5.035 1.025 5.035 1.005 5.06 1.005 5.06 0.52 4.895 0.52 4.895 0.46 5.485 0.46 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.26 0.41 9.34 0.91 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.4814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.95 0.92 8.43 0.92 8.43 0.84 8.86 0.84 8.86 0.79 8.87 0.79 8.87 0.74 8.95 0.74 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 7.26 0.78 7.39 1.23 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.54 1.04 4.46 1.04 4.46 0.73 4.4 0.73 4.4 0.65 4.46 0.65 4.46 0.6 4.54 0.6 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.59 0.985 0.19 0.985 0.19 0.805 0.58 0.805 0.58 0.905 0.59 0.905 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 17.638889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.07 0.85 1.01 0.85 1.01 0.36 0.605 0.36 0.605 0.645 0.75 0.645 0.75 0.705 0.225 0.705 0.225 0.625 0.365 0.625 0.365 0.645 0.545 0.645 0.545 0.3 1.07 0.3 ;
    END
  END SE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.6 1.77 0 1.77 0 1.65 0.385 1.65 0.385 1.245 0.505 1.245 0.505 1.305 0.445 1.305 0.445 1.65 1.245 1.65 1.245 1.54 1.365 1.54 1.365 1.65 2.105 1.65 2.105 1.51 2.165 1.51 2.165 1.65 3.505 1.65 3.505 1.54 3.625 1.54 3.625 1.65 3.89 1.65 3.89 1.54 4.01 1.54 4.01 1.65 4.5 1.65 4.5 1.49 4.62 1.49 4.62 1.55 4.56 1.55 4.56 1.65 4.97 1.65 4.97 1.49 5.09 1.49 5.09 1.55 5.03 1.55 5.03 1.65 5.47 1.65 5.47 1.49 5.59 1.49 5.59 1.55 5.53 1.55 5.53 1.65 5.94 1.65 5.94 1.46 6.06 1.46 6.06 1.52 6 1.52 6 1.65 6.41 1.65 6.41 1.49 6.53 1.49 6.53 1.55 6.47 1.55 6.47 1.65 7.305 1.65 7.305 1.51 7.365 1.51 7.365 1.65 9.155 1.65 9.155 1.34 9.275 1.34 9.275 1.4 9.215 1.4 9.215 1.65 9.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.6 0.06 9.315 0.06 9.315 0.2 9.255 0.2 9.255 0.06 8.38 0.06 8.38 0.36 8.44 0.36 8.44 0.42 8.32 0.42 8.32 0.06 8.125 0.06 8.125 0.2 8.065 0.2 8.065 0.06 7.55 0.06 7.55 0.17 7.43 0.17 7.43 0.06 6.66 0.06 6.66 0.17 6.54 0.17 6.54 0.06 6.19 0.06 6.19 0.17 6.07 0.17 6.07 0.06 5.72 0.06 5.72 0.17 5.6 0.17 5.6 0.06 5.25 0.06 5.25 0.17 5.13 0.17 5.13 0.06 4.78 0.06 4.78 0.17 4.66 0.17 4.66 0.06 3.92 0.06 3.92 0.485 3.98 0.485 3.98 0.545 3.86 0.545 3.86 0.06 3.505 0.06 3.505 0.485 3.565 0.485 3.565 0.545 3.445 0.545 3.445 0.06 2.41 0.06 2.41 0.17 2.29 0.17 2.29 0.06 1.265 0.06 1.265 0.525 1.205 0.525 1.205 0.06 0.445 0.06 0.445 0.525 0.385 0.525 0.385 0.06 0 0.06 0 -0.06 9.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 9.5 1.24 8.95 1.24 8.95 1.4 8.655 1.4 8.655 1.34 8.89 1.34 8.89 1.18 9.44 1.18 9.44 0.54 9.5 0.54 ;
      POLYGON 9.11 1.08 8.99 1.08 8.99 1.02 9.05 1.02 9.05 0.64 9.02 0.64 9.02 0.285 8.6 0.285 8.6 0.58 8.17 0.58 8.17 0.68 8.01 0.68 8.01 0.62 8.11 0.62 8.11 0.52 8.54 0.52 8.54 0.225 9.08 0.225 9.08 0.58 9.11 0.58 ;
      POLYGON 8.82 0.445 8.76 0.445 8.76 0.74 8.33 0.74 8.33 1.02 8.79 1.02 8.79 1.175 8.73 1.175 8.73 1.08 8.395 1.08 8.395 1.145 8.27 1.145 8.27 0.84 7.55 0.84 7.55 1.39 6.515 1.39 6.515 1.36 3.405 1.36 3.405 1.475 2.265 1.475 2.265 1.41 1.145 1.41 1.145 1.375 1.085 1.375 1.085 1.315 1.205 1.315 1.205 1.35 2.325 1.35 2.325 1.415 3.345 1.415 3.345 1.3 6.575 1.3 6.575 1.33 7.49 1.33 7.49 0.78 7.75 0.78 7.75 0.52 7.69 0.52 7.69 0.46 7.81 0.46 7.81 0.78 8.27 0.78 8.27 0.68 8.7 0.68 8.7 0.385 8.82 0.385 ;
      POLYGON 8.615 1.24 8.555 1.24 8.555 1.305 7.93 1.305 7.93 1.18 7.87 1.18 7.87 1.12 7.99 1.12 7.99 1.245 8.495 1.245 8.495 1.18 8.615 1.18 ;
      POLYGON 8.17 1.115 8.09 1.115 8.09 1.02 7.77 1.02 7.77 1.085 7.65 1.085 7.65 1.005 7.69 1.005 7.69 0.94 8.17 0.94 ;
      POLYGON 7.875 0.335 7.515 0.335 7.515 0.33 7.145 0.33 7.145 0.36 6.675 0.36 6.675 0.765 6.615 0.765 6.615 0.36 4.795 0.36 4.795 0.62 4.92 0.62 4.92 0.74 4.75 0.74 4.75 0.85 4.69 0.85 4.69 0.68 4.735 0.68 4.735 0.36 4.14 0.36 4.14 0.705 3.745 0.705 3.745 0.93 3.775 0.93 3.775 0.99 3.655 0.99 3.655 0.98 3.345 0.98 3.345 0.86 3.405 0.86 3.405 0.92 3.685 0.92 3.685 0.54 3.745 0.54 3.745 0.645 4.08 0.645 4.08 0.3 7.085 0.3 7.085 0.27 7.55 0.27 7.55 0.275 7.875 0.275 ;
      POLYGON 7.565 0.68 7.16 0.68 7.16 1.085 7.04 1.085 7.04 1.025 7.1 1.025 7.1 0.62 7.225 0.62 7.225 0.43 7.285 0.43 7.285 0.62 7.565 0.62 ;
      POLYGON 6.895 0.52 6.835 0.52 6.835 0.925 6.735 0.925 6.735 1.03 6.675 1.03 6.675 0.925 6.27 0.925 6.27 0.725 6.33 0.725 6.33 0.865 6.775 0.865 6.775 0.46 6.895 0.46 ;
      POLYGON 4.36 0.55 4.3 0.55 4.3 1.15 3.245 1.15 3.245 1.315 2.425 1.315 2.425 1.25 2.11 1.25 2.11 0.905 2.17 0.905 2.17 1.19 2.485 1.19 2.485 1.255 2.805 1.255 2.805 0.995 2.745 0.995 2.745 0.935 2.865 0.935 2.865 1.255 3.185 1.255 3.185 0.865 3.125 0.865 3.125 0.805 3.245 0.805 3.245 1.09 4.24 1.09 4.24 0.49 4.36 0.49 ;
      POLYGON 3.585 0.82 3.525 0.82 3.525 0.705 3.025 0.705 3.025 1.095 3.085 1.095 3.085 1.155 2.965 1.155 2.965 0.54 3.025 0.54 3.025 0.645 3.585 0.645 ;
      POLYGON 2.865 0.79 2.745 0.79 2.745 0.73 2.805 0.73 2.805 0.44 1.85 0.44 1.85 0.95 1.79 0.95 1.79 0.44 1.47 0.44 1.47 1.02 1.53 1.02 1.53 1.08 1.41 1.08 1.41 0.38 2.865 0.38 ;
      POLYGON 2.705 0.63 2.645 0.63 2.645 1.095 2.705 1.095 2.705 1.155 2.585 1.155 2.585 0.95 2.27 0.95 2.27 0.89 2.585 0.89 2.585 0.57 2.705 0.57 ;
      POLYGON 2.485 0.79 2.01 0.79 2.01 1.185 1.95 1.185 1.95 0.57 2.07 0.57 2.07 0.63 2.01 0.63 2.01 0.73 2.485 0.73 ;
      POLYGON 1.805 1.24 1.28 1.24 1.28 1.215 0.85 1.215 0.85 0.52 0.705 0.52 0.705 0.46 0.91 0.46 0.91 1.155 1.335 1.155 1.335 1.18 1.63 1.18 1.63 0.54 1.69 0.54 1.69 1.12 1.805 1.12 ;
      POLYGON 0.75 1.145 0.24 1.145 0.24 1.205 0.18 1.205 0.18 1.145 0.03 1.145 0.03 0.465 0.18 0.465 0.18 0.405 0.24 0.405 0.24 0.525 0.09 0.525 0.09 1.085 0.69 1.085 0.69 0.83 0.75 0.83 ;
  END
END SEDFFTRX4

MACRO SEDFFTRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFTRXL 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.58915 LAYER Metal1 ;
    ANTENNADIFFAREA 4.3153 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2916 LAYER Metal1 ;
      ANTENNAMAXAREACAR 15.73782575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 123.1893005 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.54 0.825 5.455 0.825 5.455 1.04 5.375 1.04 5.375 0.745 5.46 0.745 5.46 0.39 5.54 0.39 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.534725 LAYER Metal1 ;
    ANTENNADIFFAREA 4.3153 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2916 LAYER Metal1 ;
      ANTENNAMAXAREACAR 15.55118325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 122.45370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.165 0.635 0.14 0.635 0.14 1.02 0.06 1.02 0.06 0.41 0.165 0.41 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.76 1.06 7.74 1.06 7.74 1.215 7.66 1.215 7.66 0.98 7.68 0.98 7.68 0.735 7.76 0.735 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.395 0.85 7.165 0.85 7.165 0.895 7.035 0.895 7.035 0.85 6.94 0.85 6.94 0.77 7.395 0.77 ;
    END
  END E
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.07 1.015 5.94 1.015 5.94 1.25 5.86 1.25 5.86 1.015 5.805 1.015 5.805 0.935 6.07 0.935 ;
    END
  END RN
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.4074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.175 0.745 4.375 0.945 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.18518525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.755 0.705 4.695 0.705 4.695 0.645 4.075 0.645 4.075 0.705 3.835 0.705 3.835 0.625 4.015 0.625 4.015 0.585 4.755 0.585 ;
    END
  END SE
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.415 0.895 3.3 0.895 3.3 1.12 3.22 1.12 3.22 0.735 3.3 0.735 3.3 0.74 3.415 0.74 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 1.77 0 1.77 0 1.65 0.31 1.65 0.31 1.49 0.43 1.49 0.43 1.55 0.37 1.55 0.37 1.65 0.955 1.65 0.955 1.34 1.015 1.34 1.015 1.65 1.98 1.65 1.98 1.28 1.92 1.28 1.92 1.22 2.04 1.22 2.04 1.65 3.135 1.65 3.135 1.54 3.255 1.54 3.255 1.65 4.19 1.65 4.19 1.54 4.31 1.54 4.31 1.65 5.11 1.65 5.11 1.54 5.23 1.54 5.23 1.65 5.93 1.65 5.93 1.51 5.99 1.51 5.99 1.65 7.685 1.65 7.685 1.51 7.745 1.51 7.745 1.65 8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 0.06 7.715 0.06 7.715 0.635 7.655 0.635 7.655 0.06 6.925 0.06 6.925 0.29 6.985 0.29 6.985 0.35 6.865 0.35 6.865 0.06 6.64 0.06 6.64 0.29 6.7 0.29 6.7 0.35 6.58 0.35 6.58 0.06 6.145 0.06 6.145 0.515 6.025 0.515 6.025 0.455 6.085 0.455 6.085 0.06 5.2 0.06 5.2 0.485 5.14 0.485 5.14 0.06 4.25 0.06 4.25 0.265 4.31 0.265 4.31 0.325 4.19 0.325 4.19 0.06 3.195 0.06 3.195 0.475 3.135 0.475 3.135 0.06 2.04 0.06 2.04 0.28 1.92 0.28 1.92 0.22 1.98 0.22 1.98 0.06 0.985 0.06 0.985 0.635 0.925 0.635 0.925 0.06 0.37 0.06 0.37 0.635 0.31 0.635 0.31 0.06 0 0.06 0 -0.06 8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.92 1.375 7.11 1.375 7.11 1.315 7.86 1.315 7.86 0.54 7.92 0.54 ;
      POLYGON 7.555 1.01 7.51 1.01 7.51 1.07 7.45 1.07 7.45 0.95 7.495 0.95 7.495 0.67 6.625 0.67 6.625 0.73 6.565 0.73 6.565 0.61 7.42 0.61 7.42 0.57 7.54 0.57 7.54 0.61 7.555 0.61 ;
      POLYGON 7.295 0.375 7.235 0.375 7.235 0.51 6.465 0.51 6.465 0.83 6.84 0.83 6.84 0.995 7.295 0.995 7.295 1.12 7.175 1.12 7.175 1.055 6.84 1.055 6.84 1.15 6.78 1.15 6.78 0.89 6.405 0.89 6.405 0.545 6.305 0.545 6.305 0.675 5.865 0.675 5.865 0.29 5.36 0.29 5.36 0.645 5.015 0.645 5.015 0.585 5.3 0.585 5.3 0.23 5.925 0.23 5.925 0.615 6.245 0.615 6.245 0.425 6.32 0.425 6.32 0.45 7.175 0.45 7.175 0.315 7.295 0.315 ;
      POLYGON 7.075 1.215 7.01 1.215 7.01 1.355 6.4 1.355 6.4 1.29 6.375 1.29 6.375 1.17 6.435 1.17 6.435 1.235 6.46 1.235 6.46 1.295 6.95 1.295 6.95 1.155 7.075 1.155 ;
      POLYGON 6.64 1.195 6.56 1.195 6.56 1.07 6.25 1.07 6.25 1.195 6.17 1.195 6.17 0.99 6.64 0.99 ;
      POLYGON 6.3 1.425 6.18 1.425 6.18 1.41 5.01 1.41 5.01 1.44 2.14 1.44 2.14 1.12 1.82 1.12 1.82 1.375 1.235 1.375 1.235 1.44 1.115 1.44 1.115 1.24 0.54 1.24 0.54 1.245 0.42 1.245 0.42 1.185 0.48 1.185 0.48 1.18 0.69 1.18 0.69 0.57 0.81 0.57 0.81 0.63 0.75 0.63 0.75 1.18 1.175 1.18 1.175 1.315 1.76 1.315 1.76 1.06 2.2 1.06 2.2 1.38 4.95 1.38 4.95 1.35 6.24 1.35 6.24 1.365 6.3 1.365 ;
      POLYGON 6.12 0.835 5.705 0.835 5.705 1.195 5.645 1.195 5.645 0.48 5.765 0.48 5.765 0.54 5.705 0.54 5.705 0.775 6.12 0.775 ;
      POLYGON 4.925 0.225 4.64 0.225 4.64 0.485 3.735 0.485 3.735 1.045 4.475 1.045 4.475 0.79 4.595 0.79 4.595 0.85 4.535 0.85 4.535 1.105 3.675 1.105 3.675 0.425 3.985 0.425 3.985 0.365 4.045 0.365 4.045 0.425 4.58 0.425 4.58 0.165 4.925 0.165 ;
      POLYGON 4.915 1.01 4.695 1.01 4.695 1.28 2.505 1.28 2.505 1.16 2.68 1.16 2.68 0.54 2.74 0.54 2.74 1.22 4.635 1.22 4.635 0.95 4.855 0.95 4.855 0.48 4.74 0.48 4.74 0.42 4.915 0.42 ;
      POLYGON 3.575 1.055 3.4 1.055 3.4 0.995 3.515 0.995 3.515 0.635 3.12 0.635 3.12 0.695 3.06 0.695 3.06 0.575 3.515 0.575 3.515 0.475 3.37 0.475 3.37 0.355 3.43 0.355 3.43 0.415 3.575 0.415 ;
      POLYGON 2.96 1.055 2.84 1.055 2.84 0.995 2.9 0.995 2.9 0.44 2.58 0.44 2.58 1.025 2.52 1.025 2.52 0.44 1.265 0.44 1.265 0.86 1.34 0.86 1.34 0.92 1.205 0.92 1.205 0.38 1.505 0.38 1.505 0.34 1.625 0.34 1.625 0.38 2.195 0.38 2.195 0.34 2.315 0.34 2.315 0.38 2.96 0.38 ;
      POLYGON 2.42 0.63 2.36 0.63 2.36 1.215 2.3 1.215 2.3 0.8 1.815 0.8 1.815 0.74 2.3 0.74 2.3 0.57 2.42 0.57 ;
      POLYGON 2.145 0.96 1.66 0.96 1.66 1.215 1.6 1.215 1.6 0.54 1.66 0.54 1.66 0.9 2.145 0.9 ;
      POLYGON 1.5 1.215 1.395 1.215 1.395 1.08 0.86 1.08 0.86 0.91 0.92 0.91 0.92 1.02 1.44 1.02 1.44 0.63 1.365 0.63 1.365 0.57 1.5 0.57 ;
      POLYGON 0.575 1.02 0.495 1.02 0.495 0.815 0.24 0.815 0.24 0.735 0.495 0.735 0.495 0.54 0.575 0.54 ;
  END
END SEDFFTRXL

MACRO SEDFFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFX1 0 0 ;
  SIZE 7 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.7827 LAYER Metal1 ;
    ANTENNADIFFAREA 4.014875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2691 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.05685625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 111.0033445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.82 1.095 3.76 1.095 3.76 0.705 3.635 0.705 3.635 0.54 3.695 0.54 3.695 0.625 3.82 0.625 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.826 LAYER Metal1 ;
    ANTENNADIFFAREA 4.014875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2691 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.217763 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 111.8283165 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.98 0.99 1.86 0.99 1.86 0.61 1.805 0.61 1.805 0.49 1.94 0.49 1.94 0.91 1.98 0.91 ;
    END
  END QN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.66 0.79 6.88 0.98 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.62 3.34 1.12 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.445 1.06 2.34 1.06 2.34 1.12 2.26 1.12 2.26 0.98 2.365 0.98 2.365 0.725 2.445 0.725 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.54 0.815 0.88 0.935 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 23.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.52 0.91 1.46 0.91 1.46 0.395 0.945 0.395 0.945 0.655 1.04 0.655 1.04 0.78 0.98 0.78 0.98 0.715 0.44 0.715 0.44 0.895 0.235 0.895 0.235 0.815 0.38 0.815 0.38 0.655 0.885 0.655 0.885 0.335 1.52 0.335 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7 1.77 0 1.77 0 1.65 0.48 1.65 0.48 1.195 0.6 1.195 0.6 1.255 0.54 1.255 0.54 1.65 1.655 1.65 1.655 1.51 1.715 1.51 1.715 1.65 2.295 1.65 2.295 1.54 2.415 1.54 2.415 1.65 3.465 1.65 3.465 1.54 3.585 1.54 3.585 1.65 4.315 1.65 4.315 1.51 4.375 1.51 4.375 1.65 5.295 1.65 5.295 1.54 5.415 1.54 5.415 1.65 6.585 1.65 6.585 1.24 6.645 1.24 6.645 1.65 7 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7 0.06 6.56 0.06 6.56 0.53 6.5 0.53 6.5 0.06 5.425 0.06 5.425 0.16 5.485 0.16 5.485 0.22 5.365 0.22 5.365 0.06 4.44 0.06 4.44 0.215 4.5 0.215 4.5 0.275 4.38 0.275 4.38 0.06 3.375 0.06 3.375 0.52 3.315 0.52 3.315 0.06 2.315 0.06 2.315 0.625 2.255 0.625 2.255 0.06 1.545 0.06 1.545 0.2 1.485 0.2 1.485 0.06 0.545 0.06 0.545 0.555 0.425 0.555 0.425 0.495 0.485 0.495 0.485 0.06 0 0.06 0 -0.06 7 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.88 1.235 6.745 1.235 6.745 1.14 6.485 1.14 6.485 1.47 5.575 1.47 5.575 1.44 4.83 1.44 4.83 1.38 5.695 1.38 5.695 1.41 6.425 1.41 6.425 0.63 6.66 0.63 6.66 0.495 6.735 0.495 6.735 0.435 6.795 0.435 6.795 0.555 6.72 0.555 6.72 0.69 6.485 0.69 6.485 1.08 6.805 1.08 6.805 1.175 6.88 1.175 ;
      POLYGON 6.325 1.31 5.905 1.31 5.905 1.28 4.92 1.28 4.92 0.895 4.735 0.895 4.735 0.955 4.675 0.955 4.675 0.835 4.92 0.835 4.92 0.77 5.04 0.77 5.04 0.83 4.98 0.83 4.98 1.22 5.905 1.22 5.905 0.86 5.965 0.86 5.965 1.25 6.265 1.25 6.265 0.435 6.325 0.435 ;
      POLYGON 6.125 1.15 6.065 1.15 6.065 0.435 3.535 0.435 3.535 0.705 3.5 0.705 3.5 1.28 3.045 1.28 3.045 1.34 2.985 1.34 2.985 1.28 2.94 1.28 2.94 0.54 3 0.54 3 1.22 3.44 1.22 3.44 0.645 3.475 0.645 3.475 0.375 6.125 0.375 ;
      POLYGON 5.95 0.595 5.805 0.595 5.805 1.12 5.685 1.12 5.685 1.06 5.745 1.06 5.745 0.955 5.3 0.955 5.3 0.895 5.745 0.895 5.745 0.535 5.95 0.535 ;
      POLYGON 5.56 0.795 5.5 0.795 5.5 0.735 5.2 0.735 5.2 1.12 5.08 1.12 5.08 1.06 5.14 1.06 5.14 0.595 4.985 0.595 4.985 0.535 5.2 0.535 5.2 0.675 5.56 0.675 ;
      POLYGON 4.885 0.595 4.82 0.595 4.82 0.735 4.575 0.735 4.575 1.06 4.82 1.06 4.82 1.12 4.515 1.12 4.515 0.915 4.19 0.915 4.19 0.855 4.515 0.855 4.515 0.675 4.76 0.675 4.76 0.535 4.885 0.535 ;
      POLYGON 4.415 0.755 4.06 0.755 4.06 1.015 4.14 1.015 4.14 1.44 3.205 1.44 3.205 1.5 2.515 1.5 2.515 1.44 2.135 1.44 2.135 1.38 2.575 1.38 2.575 1.44 3.145 1.44 3.145 1.38 3.6 1.38 3.6 0.805 3.66 0.805 3.66 1.38 4.08 1.38 4.08 1.075 4 1.075 4 0.535 4.12 0.535 4.12 0.595 4.06 0.595 4.06 0.695 4.415 0.695 ;
      POLYGON 3.16 1.055 3.1 1.055 3.1 0.255 2.52 0.255 2.52 0.565 2.605 0.565 2.605 0.73 2.62 0.73 2.62 1.08 2.56 1.08 2.56 0.79 2.545 0.79 2.545 0.625 2.46 0.625 2.46 0.195 3.16 0.195 ;
      POLYGON 2.84 1.28 1.3 1.28 1.3 0.555 1.045 0.555 1.045 0.495 1.36 0.495 1.36 1.22 2.765 1.22 2.765 0.63 2.705 0.63 2.705 0.57 2.825 0.57 2.825 1.16 2.84 1.16 ;
      POLYGON 2.15 1.08 2.09 1.08 2.09 0.625 2.05 0.625 2.05 0.39 1.705 0.39 1.705 0.795 1.645 0.795 1.645 0.33 2.11 0.33 2.11 0.565 2.15 0.565 ;
      POLYGON 1.2 1.095 0.365 1.095 0.365 1.19 0.305 1.19 0.305 1.095 0.075 1.095 0.075 0.55 0.22 0.55 0.22 0.49 0.28 0.49 0.28 0.61 0.135 0.61 0.135 1.035 1.14 1.035 1.14 0.91 1.2 0.91 ;
  END
END SEDFFX1

MACRO SEDFFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFX2 0 0 ;
  SIZE 7.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.332675 LAYER Metal1 ;
    ANTENNADIFFAREA 4.2666 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.334575 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.949787 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 101.241874 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.18 1.11 6.06 1.11 6.06 0.98 6.1 0.98 6.1 0.4 6.18 0.4 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.285075 LAYER Metal1 ;
    ANTENNADIFFAREA 4.2666 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.334575 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.807517 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 100.49764625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.34 1.29 0.28 1.29 0.28 0.73 0.26 0.73 0.26 0.6 0.28 0.6 0.28 0.54 0.34 0.54 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.425926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.565 0.705 7.425 0.705 7.425 0.645 6.795 0.645 6.795 0.65 6.735 0.65 6.735 1.085 6.675 1.085 6.675 0.585 7.485 0.585 7.485 0.625 7.565 0.625 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.325 0.825 7.165 0.825 7.165 0.895 6.895 0.895 6.895 0.745 7.325 0.745 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.62962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.635 0.61 5.765 0.98 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.365 1.265 4.285 1.265 4.285 0.895 4.235 0.895 4.235 0.815 4.365 0.815 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.135 1.06 4.055 1.06 4.055 0.92 3.86 0.92 3.86 0.755 3.94 0.755 3.94 0.84 4.135 0.84 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.8 1.77 0 1.77 0 1.65 0.075 1.65 0.075 0.9 0.135 0.9 0.135 1.65 0.515 1.65 0.515 1.51 0.575 1.51 0.575 1.65 0.87 1.65 0.87 1.35 0.93 1.35 0.93 1.65 1.905 1.65 1.905 1.28 1.845 1.28 1.845 1.22 1.965 1.22 1.965 1.65 3.06 1.65 3.06 1.31 3 1.31 3 1.25 3.12 1.25 3.12 1.65 4.205 1.65 4.205 1.54 4.325 1.54 4.325 1.65 5.825 1.65 5.825 1.42 5.945 1.42 5.945 1.48 5.885 1.48 5.885 1.65 6.295 1.65 6.295 1.42 6.415 1.42 6.415 1.48 6.355 1.48 6.355 1.65 7.11 1.65 7.11 1.22 7.17 1.22 7.17 1.65 7.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.8 0.06 7.065 0.06 7.065 0.405 7.125 0.405 7.125 0.465 7.005 0.465 7.005 0.06 6.395 0.06 6.395 0.2 6.335 0.2 6.335 0.06 5.985 0.06 5.985 0.35 5.865 0.35 5.865 0.29 5.925 0.29 5.925 0.06 4.395 0.06 4.395 0.495 4.335 0.495 4.335 0.06 3.185 0.06 3.185 0.635 3.125 0.635 3.125 0.06 1.965 0.06 1.965 0.28 1.845 0.28 1.845 0.22 1.905 0.22 1.905 0.06 1.03 0.06 1.03 0.2 0.97 0.2 0.97 0.06 0.545 0.06 0.545 0.52 0.485 0.52 0.485 0.06 0.135 0.06 0.135 0.52 0.075 0.52 0.075 0.06 0 0.06 0 -0.06 7.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.725 1.215 7.56 1.215 7.56 1.275 7.5 1.275 7.5 1.155 7.665 1.155 7.665 1.055 6.835 1.055 6.835 0.995 7.665 0.995 7.665 0.485 7.47 0.485 7.47 0.425 7.725 0.425 ;
      POLYGON 6.83 1.32 4.9 1.32 4.9 1.095 5.09 1.095 5.09 0.49 4.975 0.49 4.975 0.43 5.15 0.43 5.15 1.155 4.96 1.155 4.96 1.26 6.515 1.26 6.515 0.425 6.755 0.425 6.755 0.485 6.575 0.485 6.575 1.25 6.83 1.25 ;
      POLYGON 6 0.88 5.94 0.88 5.94 0.51 5.705 0.51 5.705 0.33 4.555 0.33 4.555 0.655 4.175 0.655 4.175 0.33 3.39 0.33 3.39 0.635 3.6 0.635 3.6 1.02 3.54 1.02 3.54 0.695 3.33 0.695 3.33 0.27 4.235 0.27 4.235 0.595 4.495 0.595 4.495 0.27 5.765 0.27 5.765 0.45 6 0.45 ;
      POLYGON 5.635 1.16 5.25 1.16 5.25 0.43 5.605 0.43 5.605 0.51 5.33 0.51 5.33 0.61 5.37 0.61 5.37 0.69 5.33 0.69 5.33 1.08 5.635 1.08 ;
      POLYGON 4.99 0.995 4.625 0.995 4.625 0.915 4.91 0.915 4.91 0.595 4.99 0.595 ;
      POLYGON 4.81 0.49 4.715 0.49 4.715 0.815 4.525 0.815 4.525 1.095 4.705 1.095 4.705 1.215 4.645 1.215 4.645 1.155 4.525 1.155 4.525 1.44 3.22 1.44 3.22 1.15 2.52 1.15 2.52 1.215 2.46 1.215 2.46 1.09 2.605 1.09 2.605 0.54 2.665 0.54 2.665 1.09 3.28 1.09 3.28 1.38 4.465 1.38 4.465 0.755 4.655 0.755 4.655 0.43 4.81 0.43 ;
      POLYGON 4.075 0.49 3.76 0.49 3.76 1.16 4.06 1.16 4.06 1.28 4 1.28 4 1.22 3.38 1.22 3.38 0.855 2.985 0.855 2.985 0.735 3.045 0.735 3.045 0.795 3.44 0.795 3.44 1.16 3.7 1.16 3.7 0.43 4.075 0.43 ;
      POLYGON 2.98 0.635 2.885 0.635 2.885 0.99 2.765 0.99 2.765 0.93 2.825 0.93 2.825 0.575 2.92 0.575 2.92 0.475 2.765 0.475 2.765 0.44 2.505 0.44 2.505 0.91 2.445 0.91 2.445 0.97 2.385 0.97 2.385 0.85 2.445 0.85 2.445 0.44 1.685 0.44 1.685 0.4 1.19 0.4 1.19 0.87 1.265 0.87 1.265 0.93 1.13 0.93 1.13 0.34 1.745 0.34 1.745 0.38 2.12 0.38 2.12 0.34 2.24 0.34 2.24 0.38 2.825 0.38 2.825 0.415 2.98 0.415 ;
      POLYGON 2.9 1.405 2.065 1.405 2.065 1.12 1.745 1.12 1.745 1.375 1.15 1.375 1.15 1.44 1.03 1.44 1.03 1.38 1.09 1.38 1.09 1.25 0.715 1.25 0.715 0.99 0.645 0.99 0.645 0.79 0.44 0.79 0.44 0.73 0.645 0.73 0.645 0.57 0.81 0.57 0.81 0.63 0.705 0.63 0.705 0.93 0.775 0.93 0.775 1.19 1.15 1.19 1.15 1.315 1.685 1.315 1.685 1.06 2.125 1.06 2.125 1.345 2.9 1.345 ;
      POLYGON 2.345 0.63 2.285 0.63 2.285 1.215 2.225 1.215 2.225 0.8 1.74 0.8 1.74 0.74 2.225 0.74 2.225 0.57 2.345 0.57 ;
      POLYGON 2.06 0.96 1.585 0.96 1.585 1.215 1.525 1.215 1.525 0.54 1.585 0.54 1.585 0.9 2.06 0.9 ;
      POLYGON 1.425 1.185 1.29 1.185 1.29 1.09 0.97 1.09 0.97 0.83 0.805 0.83 0.805 0.77 1.03 0.77 1.03 1.03 1.365 1.03 1.365 0.63 1.29 0.63 1.29 0.57 1.425 0.57 ;
  END
END SEDFFX2

MACRO SEDFFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFX4 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5419 LAYER Metal1 ;
    ANTENNADIFFAREA 4.865175 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4878 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.310988 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 73.198032 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.675 0.625 6.32 0.625 6.32 0.98 6.34 0.98 6.34 1.005 6.575 1.005 6.575 1.02 6.635 1.02 6.635 1.08 6.515 1.08 6.515 1.065 6.34 1.065 6.34 1.11 6.045 1.11 6.045 1.05 6.26 1.05 6.26 0.625 6.205 0.625 6.205 0.485 6.265 0.485 6.265 0.565 6.615 0.565 6.615 0.485 6.675 0.485 ;
    END
  END QN
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 9.72222225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.74 0.785 7.35 0.785 7.35 0.855 7.105 0.855 7.105 0.955 7.045 0.955 7.045 0.795 7.29 0.795 7.29 0.725 7.46 0.725 7.46 0.6 7.54 0.6 7.54 0.725 7.74 0.725 ;
    END
  END E
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.795 1.085 7.54 1.085 7.54 1.11 7.44 1.11 7.44 0.98 7.45 0.98 7.45 0.885 7.795 0.885 ;
    END
  END D
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.94 0.925 5.91 0.925 5.91 1.195 5.83 1.195 5.83 0.725 5.94 0.725 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.765 0.96 4.685 0.96 4.685 0.59 4.635 0.59 4.635 0.51 4.765 0.51 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.962963 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.435 0.69 4.575 0.98 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5419 LAYER Metal1 ;
    ANTENNADIFFAREA 4.865175 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4878 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.310988 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 73.198032 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.745 0.66 0.7 0.66 0.7 0.915 0.745 0.915 0.745 1.345 0.685 1.345 0.685 0.975 0.64 0.975 0.64 0.73 0.335 0.73 0.335 1.345 0.26 1.345 0.26 0.54 0.335 0.54 0.335 0.6 0.34 0.6 0.34 0.67 0.64 0.67 0.64 0.6 0.685 0.6 0.685 0.54 0.745 0.54 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 1.77 0 1.77 0 1.65 0.07 1.65 0.07 0.955 0.13 0.955 0.13 1.65 0.48 1.65 0.48 0.955 0.54 0.955 0.54 1.65 0.89 1.65 0.89 1.035 0.95 1.035 0.95 1.65 1.33 1.65 1.33 1.32 1.39 1.32 1.39 1.65 2.385 1.65 2.385 1.22 2.325 1.22 2.325 1.16 2.445 1.16 2.445 1.65 3.56 1.65 3.56 1.31 3.5 1.31 3.5 1.25 3.62 1.25 3.62 1.65 4.64 1.65 4.64 1.24 4.7 1.24 4.7 1.65 5.81 1.65 5.81 1.455 5.93 1.455 5.93 1.515 5.87 1.515 5.87 1.65 6.28 1.65 6.28 1.455 6.4 1.455 6.4 1.515 6.34 1.515 6.34 1.65 6.75 1.65 6.75 1.455 6.87 1.455 6.87 1.515 6.81 1.515 6.81 1.65 7.555 1.65 7.555 1.51 7.615 1.51 7.615 1.65 8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 0.06 7.64 0.06 7.64 0.5 7.58 0.5 7.58 0.06 6.88 0.06 6.88 0.465 6.82 0.465 6.82 0.06 6.47 0.06 6.47 0.465 6.41 0.465 6.41 0.06 6.06 0.06 6.06 0.465 6 0.465 6 0.06 4.715 0.06 4.715 0.25 4.595 0.25 4.595 0.19 4.655 0.19 4.655 0.06 3.665 0.06 3.665 0.52 3.605 0.52 3.605 0.06 2.445 0.06 2.445 0.25 2.325 0.25 2.325 0.19 2.385 0.19 2.385 0.06 1.39 0.06 1.39 0.575 1.33 0.575 1.33 0.06 0.95 0.06 0.95 0.52 0.89 0.52 0.89 0.06 0.54 0.06 0.54 0.52 0.48 0.52 0.48 0.06 0.13 0.06 0.13 0.52 0.07 0.52 0.07 0.06 0 0.06 0 -0.06 8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.955 1.33 7.79 1.33 7.79 1.27 7.28 1.27 7.28 0.955 7.34 0.955 7.34 1.21 7.895 1.21 7.895 0.525 7.785 0.525 7.785 0.405 7.845 0.405 7.845 0.465 7.955 0.465 ;
      POLYGON 7.255 0.625 6.945 0.625 6.945 1.21 7.18 1.21 7.18 1.355 5.3 1.355 5.3 0.91 5.49 0.91 5.49 0.59 5.405 0.59 5.405 0.47 5.465 0.47 5.465 0.53 5.55 0.53 5.55 0.97 5.36 0.97 5.36 1.295 6.885 1.295 6.885 0.565 7.195 0.565 7.195 0.405 7.255 0.405 ;
      POLYGON 6.105 0.765 6.045 0.765 6.045 0.625 5.84 0.625 5.84 0.385 5.565 0.385 5.565 0.37 5.05 0.37 5.05 0.41 4.435 0.41 4.435 0.37 3.87 0.37 3.87 0.47 4.1 0.47 4.1 1.02 4.04 1.02 4.04 0.53 3.81 0.53 3.81 0.31 4.495 0.31 4.495 0.35 4.99 0.35 4.99 0.31 5.625 0.31 5.625 0.325 5.9 0.325 5.9 0.565 6.105 0.565 ;
      POLYGON 5.74 0.605 5.73 0.605 5.73 1.15 5.575 1.15 5.575 1.07 5.65 1.07 5.65 0.525 5.66 0.525 5.66 0.485 5.74 0.485 ;
      POLYGON 5.39 0.81 5.145 0.81 5.145 1.05 5.025 1.05 5.025 0.97 5.065 0.97 5.065 0.73 5.31 0.73 5.31 0.69 5.39 0.69 ;
      POLYGON 5.21 0.615 4.925 0.615 4.925 1.175 5.125 1.175 5.125 1.235 4.865 1.235 4.865 1.14 4.54 1.14 4.54 1.425 3.72 1.425 3.72 1.15 2.97 1.15 2.97 1.21 2.91 1.21 2.91 1.09 3.085 1.09 3.085 0.48 3.145 0.48 3.145 1.09 3.78 1.09 3.78 1.365 4.48 1.365 4.48 1.08 4.865 1.08 4.865 0.555 5.15 0.555 5.15 0.495 5.21 0.495 ;
      POLYGON 4.38 1.265 3.88 1.265 3.88 0.815 3.405 0.815 3.405 0.755 3.94 0.755 3.94 1.205 4.275 1.205 4.275 0.47 4.335 0.47 4.335 1.145 4.38 1.145 ;
      POLYGON 3.43 0.655 3.305 0.655 3.305 0.93 3.385 0.93 3.385 0.99 3.245 0.99 3.245 0.595 3.37 0.595 3.37 0.495 3.245 0.495 3.245 0.38 2.985 0.38 2.985 0.92 2.865 0.92 2.865 0.86 2.925 0.86 2.925 0.38 2.605 0.38 2.605 0.41 2.165 0.41 2.165 0.38 1.67 0.38 1.67 0.9 1.61 0.9 1.61 0.32 1.91 0.32 1.91 0.28 2.03 0.28 2.03 0.32 2.225 0.32 2.225 0.35 2.545 0.35 2.545 0.32 2.6 0.32 2.6 0.28 2.72 0.28 2.72 0.32 3.305 0.32 3.305 0.435 3.43 0.435 ;
      POLYGON 3.4 1.405 2.545 1.405 2.545 1.06 2.225 1.06 2.225 1.315 1.61 1.315 1.61 1.38 1.49 1.38 1.49 1.22 1.155 1.22 1.155 1.345 1.095 1.345 1.095 1.095 1.05 1.095 1.05 0.815 0.8 0.815 0.8 0.755 1.05 0.755 1.05 0.72 1.125 0.72 1.125 0.54 1.185 0.54 1.185 0.78 1.11 0.78 1.11 1.035 1.155 1.035 1.155 1.16 1.55 1.16 1.55 1.255 2.165 1.255 2.165 1 2.605 1 2.605 1.345 3.4 1.345 ;
      POLYGON 2.825 0.57 2.765 0.57 2.765 1.155 2.705 1.155 2.705 0.74 2.22 0.74 2.22 0.68 2.705 0.68 2.705 0.51 2.825 0.51 ;
      POLYGON 2.55 0.9 2.065 0.9 2.065 1.155 2.005 1.155 2.005 0.48 2.065 0.48 2.065 0.84 2.55 0.84 ;
      POLYGON 1.89 0.57 1.83 0.57 1.83 1.065 1.89 1.065 1.89 1.125 1.77 1.125 1.77 1.06 1.27 1.06 1.27 0.94 1.21 0.94 1.21 0.88 1.33 0.88 1.33 1 1.77 1 1.77 0.51 1.89 0.51 ;
  END
END SEDFFX4

MACRO SEDFFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SEDFFXL 0 0 ;
  SIZE 7.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.9285 LAYER Metal1 ;
    ANTENNADIFFAREA 3.899675 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.243 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.16666675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 126.580247 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.98 1.16 3.86 1.16 3.86 0.5 3.845 0.5 3.845 0.375 3.925 0.375 3.925 0.42 3.94 0.42 3.94 1.08 3.98 1.08 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.8649 LAYER Metal1 ;
    ANTENNADIFFAREA 3.899675 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.243 LAYER Metal1 ;
      ANTENNAMAXAREACAR 15.90493825 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 125.5 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.775 1.21 1.695 1.21 1.695 0.73 1.66 0.73 1.66 0.68 1.63 0.68 1.63 0.48 1.71 0.48 1.71 0.6 1.74 0.6 1.74 0.65 1.775 0.65 ;
    END
  END QN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.17 0.91 6.94 0.91 6.94 1.06 6.86 1.06 6.86 0.79 7.17 0.79 ;
    END
  END CK
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.46 0.57 3.54 1.07 ;
    END
  END SI
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.52 0.895 2.34 0.895 2.34 0.975 2.26 0.975 2.26 0.735 2.34 0.735 2.34 0.815 2.44 0.815 2.44 0.735 2.52 0.735 ;
    END
  END SE
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.77777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.805 0.705 0.955 ;
    END
  END D
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 20.60185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.345 0.93 1.285 0.93 1.285 0.385 0.765 0.385 0.765 0.645 0.865 0.645 0.865 0.77 0.805 0.77 0.805 0.705 0.335 0.705 0.335 0.77 0.275 0.77 0.275 0.645 0.635 0.645 0.635 0.625 0.705 0.625 0.705 0.325 1.345 0.325 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 1.77 0 1.77 0 1.65 0.51 1.65 0.51 1.215 0.63 1.215 0.63 1.275 0.57 1.275 0.57 1.65 1.55 1.65 1.55 1.51 1.61 1.51 1.61 1.65 2.385 1.65 2.385 1.54 2.505 1.54 2.505 1.65 3.525 1.65 3.525 1.49 3.645 1.49 3.645 1.55 3.585 1.55 3.585 1.65 4.43 1.65 4.43 1.055 4.49 1.055 4.49 1.65 5.515 1.65 5.515 1.54 5.635 1.54 5.635 1.65 6.725 1.65 6.725 1.415 6.845 1.415 6.845 1.475 6.785 1.475 6.785 1.65 7.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 0.06 6.815 0.06 6.815 0.53 6.755 0.53 6.755 0.06 5.69 0.06 5.69 0.25 5.57 0.25 5.57 0.19 5.63 0.19 5.63 0.06 4.6 0.06 4.6 0.25 4.48 0.25 4.48 0.19 4.54 0.19 4.54 0.06 3.585 0.06 3.585 0.47 3.525 0.47 3.525 0.06 2.445 0.06 2.445 0.635 2.385 0.635 2.385 0.06 1.37 0.06 1.37 0.2 1.31 0.2 1.31 0.06 0.44 0.06 0.44 0.545 0.38 0.545 0.38 0.06 0 0.06 0 -0.06 7.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.08 1.22 6.74 1.22 6.74 1.315 6.625 1.315 6.625 1.4 4.935 1.4 4.935 1.31 5.055 1.31 5.055 1.34 6.565 1.34 6.565 1.255 6.68 1.255 6.68 0.63 6.915 0.63 6.915 0.495 6.99 0.495 6.99 0.435 7.05 0.435 7.05 0.555 6.975 0.555 6.975 0.69 6.74 0.69 6.74 1.16 7.08 1.16 ;
      POLYGON 6.58 1.155 6.465 1.155 6.465 1.24 6.085 1.24 6.085 1.21 5.105 1.21 5.105 0.89 4.82 0.89 4.82 0.83 5.225 0.83 5.225 0.89 5.165 0.89 5.165 1.15 6.085 1.15 6.085 0.89 6.025 0.89 6.025 0.83 6.145 0.83 6.145 1.18 6.405 1.18 6.405 1.095 6.52 1.095 6.52 0.435 6.58 0.435 ;
      POLYGON 6.305 1.08 6.245 1.08 6.245 0.41 4.32 0.41 4.32 0.275 3.745 0.275 3.745 1.23 3.08 1.23 3.08 0.405 3.2 0.405 3.2 0.465 3.14 0.465 3.14 1.17 3.685 1.17 3.685 0.215 4.38 0.215 4.38 0.35 6.305 0.35 ;
      POLYGON 6.13 0.57 5.925 0.57 5.925 0.99 5.985 0.99 5.985 1.05 5.865 1.05 5.865 0.93 5.545 0.93 5.545 0.865 5.485 0.865 5.485 0.805 5.605 0.805 5.605 0.87 5.865 0.87 5.865 0.51 6.13 0.51 ;
      POLYGON 5.765 0.77 5.705 0.77 5.705 0.705 5.385 0.705 5.385 1.05 5.265 1.05 5.265 0.99 5.325 0.99 5.325 0.57 5.19 0.57 5.19 0.51 5.385 0.51 5.385 0.645 5.765 0.645 ;
      POLYGON 5.085 0.57 4.72 0.57 4.72 0.99 4.895 0.99 4.895 1.05 4.66 1.05 4.66 0.89 4.26 0.89 4.26 0.83 4.66 0.83 4.66 0.51 5.085 0.51 ;
      POLYGON 4.56 0.73 4.16 0.73 4.16 0.99 4.285 0.99 4.285 1.39 2.605 1.39 2.605 1.325 2.225 1.325 2.225 1.265 2.665 1.265 2.665 1.33 4.225 1.33 4.225 1.05 4.1 1.05 4.1 0.51 4.22 0.51 4.22 0.57 4.16 0.57 4.16 0.67 4.56 0.67 ;
      POLYGON 3.36 0.855 3.24 0.855 3.24 0.795 3.3 0.795 3.3 0.305 2.65 0.305 2.65 0.595 2.68 0.595 2.68 0.945 2.74 0.945 2.74 1.005 2.62 1.005 2.62 0.655 2.59 0.655 2.59 0.245 2.99 0.245 2.99 0.17 3.11 0.17 3.11 0.245 3.36 0.245 ;
      POLYGON 2.98 1.165 2.125 1.165 2.125 1.37 1.125 1.37 1.125 0.545 0.865 0.545 0.865 0.485 1.185 0.485 1.185 1.31 2.065 1.31 2.065 1.105 2.92 1.105 2.92 0.465 2.86 0.465 2.86 0.405 2.98 0.405 ;
      POLYGON 2.16 1.005 2.04 1.005 2.04 0.945 2.1 0.945 2.1 0.5 1.81 0.5 1.81 0.38 1.53 0.38 1.53 0.785 1.47 0.785 1.47 0.32 1.87 0.32 1.87 0.44 2.16 0.44 ;
      POLYGON 1.025 1.115 0.395 1.115 0.395 1.21 0.335 1.21 0.335 1.115 0.115 1.115 0.115 0.515 0.135 0.515 0.135 0.455 0.195 0.455 0.195 0.575 0.175 0.575 0.175 1.055 0.965 1.055 0.965 0.92 1.025 0.92 ;
  END
END SEDFFXL

MACRO SMDFFHQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SMDFFHQX1 0 0 ;
  SIZE 6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1695 LAYER Metal1 ;
    ANTENNADIFFAREA 3.849 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.28935 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.953862 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 86.93105225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.145 1.34 0.085 1.34 0.085 0.73 0.06 0.73 0.06 0.6 0.085 0.6 0.085 0.54 0.145 0.54 ;
    END
  END Q
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.349835 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.79 0.765 5.73 0.765 5.73 0.705 5.135 0.705 5.135 0.83 5.06 0.83 5.06 1.04 5 1.04 5 0.77 5.075 0.77 5.075 0.645 5.235 0.645 5.235 0.625 5.365 0.625 5.365 0.645 5.79 0.645 ;
    END
  END S0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.63 1.085 5.55 1.085 5.55 0.925 5.33 0.925 5.33 0.805 5.63 0.805 ;
    END
  END D1
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.66 0.485 4.74 0.985 ;
    END
  END D0
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.82838275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.46 0.6 4.54 1.1 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.615 1.01 3.535 1.01 3.535 0.82 3.46 0.82 3.46 0.585 3.54 0.585 3.54 0.6 3.615 0.6 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.51 1 0.34 1 0.34 1.11 0.26 1.11 0.26 0.92 0.43 0.92 0.43 0.78 0.51 0.78 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 1.77 0 1.77 0 1.65 0.29 1.65 0.29 1.22 0.35 1.22 0.35 1.65 1.215 1.65 1.215 1.315 1.335 1.315 1.335 1.375 1.275 1.375 1.275 1.65 2.41 1.65 2.41 1.315 2.53 1.315 2.53 1.375 2.47 1.375 2.47 1.65 3.525 1.65 3.525 1.27 3.585 1.27 3.585 1.65 4.7 1.65 4.7 1.36 4.76 1.36 4.76 1.65 5.52 1.65 5.52 1.36 5.58 1.36 5.58 1.65 6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 0.06 5.58 0.06 5.58 0.5 5.52 0.5 5.52 0.06 4.795 0.06 4.795 0.385 4.735 0.385 4.735 0.06 3.73 0.06 3.73 0.485 3.67 0.485 3.67 0.06 2.53 0.06 2.53 0.17 2.41 0.17 2.41 0.06 1.19 0.06 1.19 0.345 1.25 0.345 1.25 0.405 1.13 0.405 1.13 0.06 0.35 0.06 0.35 0.52 0.29 0.52 0.29 0.06 0 0.06 0 -0.06 6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.95 1.245 5.815 1.245 5.815 1.305 5.755 1.305 5.755 1.245 5.17 1.245 5.17 0.93 5.23 0.93 5.23 1.185 5.89 1.185 5.89 0.525 5.755 0.525 5.755 0.405 5.815 0.405 5.815 0.465 5.95 0.465 ;
      POLYGON 5.27 0.44 4.975 0.44 4.975 0.67 4.9 0.67 4.9 1.2 5.07 1.2 5.07 1.48 5.01 1.48 5.01 1.26 4.225 1.26 4.225 1.14 4.3 1.14 4.3 0.505 4.36 0.505 4.36 1.2 4.84 1.2 4.84 0.61 4.915 0.61 4.915 0.38 5.21 0.38 5.21 0.32 5.27 0.32 ;
      POLYGON 4.56 0.5 4.5 0.5 4.5 0.405 4.2 0.405 4.2 0.95 4.125 0.95 4.125 1.36 4.555 1.36 4.555 1.48 4.495 1.48 4.495 1.42 4.065 1.42 4.065 0.95 3.875 0.95 3.875 0.83 3.935 0.83 3.935 0.89 4.14 0.89 4.14 0.345 4.56 0.345 ;
      POLYGON 4.04 0.73 3.775 0.73 3.775 1.11 3.965 1.11 3.965 1.39 3.905 1.39 3.905 1.17 3.295 1.17 3.295 1.055 3.235 1.055 3.235 0.995 3.295 0.995 3.295 0.49 3.235 0.49 3.235 0.43 3.355 0.43 3.355 1.11 3.715 1.11 3.715 0.67 3.98 0.67 3.98 0.505 4.04 0.505 ;
      POLYGON 3.525 0.485 3.465 0.485 3.465 0.33 3.135 0.33 3.135 1.27 3.41 1.27 3.41 1.33 3.075 1.33 3.075 0.33 2.755 0.33 2.755 0.625 2.815 0.625 2.815 0.685 2.695 0.685 2.695 0.33 1.93 0.33 1.93 0.59 2.045 0.59 2.045 0.71 1.985 0.71 1.985 0.65 1.87 0.65 1.87 0.27 3.525 0.27 ;
      POLYGON 2.975 1.245 2.915 1.245 2.915 0.845 2.305 0.845 2.305 0.785 2.915 0.785 2.915 0.49 2.855 0.49 2.855 0.43 2.975 0.43 ;
      POLYGON 2.865 1.405 2.745 1.405 2.745 1.215 1.885 1.215 1.885 1.26 1.435 1.26 1.435 1.215 0.61 1.215 0.61 0.54 0.67 0.54 0.67 1.155 1.435 1.155 1.435 0.725 1.385 0.725 1.385 0.665 1.505 0.665 1.505 0.725 1.495 0.725 1.495 1.2 1.825 1.2 1.825 0.88 1.765 0.88 1.765 0.82 1.885 0.82 1.885 1.155 2.805 1.155 2.805 1.345 2.865 1.345 ;
      POLYGON 2.595 0.65 2.205 0.65 2.205 1.055 2.085 1.055 2.085 0.995 2.145 0.995 2.145 0.49 2.03 0.49 2.03 0.43 2.205 0.43 2.205 0.59 2.595 0.59 ;
      POLYGON 1.725 1.1 1.665 1.1 1.665 1.04 1.605 1.04 1.605 0.565 1.145 0.565 1.145 0.69 1.085 0.69 1.085 0.505 1.605 0.505 1.605 0.4 1.665 0.4 1.665 0.98 1.725 0.98 ;
      POLYGON 1.335 0.885 0.985 0.885 0.985 0.995 1.1 0.995 1.1 1.055 0.925 1.055 0.925 0.44 0.51 0.44 0.51 0.68 0.305 0.68 0.305 0.82 0.245 0.82 0.245 0.62 0.45 0.62 0.45 0.38 0.985 0.38 0.985 0.825 1.335 0.825 ;
  END
END SMDFFHQX1

MACRO SMDFFHQX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SMDFFHQX2 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.4287 LAYER Metal1 ;
    ANTENNADIFFAREA 4.187275 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.324675 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.5604065 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 83.19242325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.355 1.31 0.295 1.31 0.295 0.92 0.26 0.92 0.26 0.79 0.28 0.79 0.28 0.54 0.34 0.54 0.34 0.875 0.355 0.875 ;
    END
  END Q
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.4158415 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.315 0.745 6.255 0.745 6.255 0.705 5.735 0.705 5.735 0.755 5.52 0.755 5.52 0.945 5.4 0.945 5.4 0.885 5.46 0.885 5.46 0.695 5.675 0.695 5.675 0.645 6.035 0.645 6.035 0.625 6.315 0.625 ;
    END
  END S0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.155 1.01 5.78 1.01 5.78 0.885 5.835 0.885 5.835 0.805 6.155 0.805 ;
    END
  END D1
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.14 0.93 4.945 0.93 4.945 0.85 5.06 0.85 5.06 0.545 5.14 0.545 ;
    END
  END D0
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.82838275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.94 0.73 4.845 0.73 4.845 0.945 4.765 0.945 4.765 0.65 4.86 0.65 4.86 0.54 4.94 0.54 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.92 0.92 3.66 0.92 3.66 0.79 3.74 0.79 3.74 0.84 3.84 0.84 3.84 0.65 3.92 0.65 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.75 0.74 1.25 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 1.77 0 1.77 0 1.65 0.09 1.65 0.09 0.92 0.15 0.92 0.15 1.65 0.5 1.65 0.5 0.92 0.56 0.92 0.56 1.65 1.33 1.65 1.33 1.25 1.45 1.25 1.45 1.31 1.39 1.31 1.39 1.65 2.61 1.65 2.61 1.405 2.73 1.405 2.73 1.465 2.67 1.465 2.67 1.65 3.82 1.65 3.82 1.225 3.88 1.225 3.88 1.65 5.15 1.65 5.15 1.205 5.21 1.205 5.21 1.65 5.885 1.65 5.885 1.285 5.945 1.285 5.945 1.65 6.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 0.06 6.02 0.06 6.02 0.525 5.96 0.525 5.96 0.06 5.21 0.06 5.21 0.435 5.15 0.435 5.15 0.06 3.95 0.06 3.95 0.545 3.89 0.545 3.89 0.06 2.795 0.06 2.795 0.475 2.675 0.475 2.675 0.415 2.735 0.415 2.735 0.06 1.47 0.06 1.47 0.49 1.35 0.49 1.35 0.43 1.41 0.43 1.41 0.06 0.515 0.06 0.515 0.43 0.575 0.43 0.575 0.49 0.455 0.49 0.455 0.06 0.135 0.06 0.135 0.52 0.075 0.52 0.075 0.06 0 0.06 0 -0.06 6.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.475 1.17 6.18 1.17 6.18 1.23 6.12 1.23 6.12 1.17 5.62 1.17 5.62 0.855 5.68 0.855 5.68 1.11 6.415 1.11 6.415 0.43 6.475 0.43 ;
      POLYGON 5.71 0.545 5.37 0.545 5.37 0.595 5.3 0.595 5.3 1.045 5.52 1.045 5.52 1.405 5.46 1.405 5.46 1.105 4.51 1.105 4.51 1.165 4.45 1.165 4.45 1.045 4.605 1.045 4.605 0.465 4.725 0.465 4.725 0.525 4.665 0.525 4.665 1.045 5.24 1.045 5.24 0.535 5.31 0.535 5.31 0.485 5.65 0.485 5.65 0.425 5.71 0.425 ;
      POLYGON 5.005 1.325 4.29 1.325 4.29 0.905 4.18 0.905 4.18 0.785 4.24 0.785 4.24 0.845 4.445 0.845 4.445 0.305 4.895 0.305 4.895 0.44 4.835 0.44 4.835 0.365 4.505 0.365 4.505 0.905 4.35 0.905 4.35 1.265 4.945 1.265 4.945 1.205 5.005 1.205 ;
      POLYGON 4.345 0.575 4.11 0.575 4.11 0.685 4.08 0.685 4.08 1.02 4.19 1.02 4.19 1.345 4.13 1.345 4.13 1.08 3.515 1.08 3.515 1.145 3.455 1.145 3.455 0.515 3.575 0.515 3.575 0.575 3.515 0.575 3.515 1.02 4.02 1.02 4.02 0.625 4.05 0.625 4.05 0.515 4.345 0.515 ;
      POLYGON 3.745 0.545 3.685 0.545 3.685 0.415 3.355 0.415 3.355 1.255 3.705 1.255 3.705 1.315 3.295 1.315 3.295 0.415 2.975 0.415 2.975 0.675 3.035 0.675 3.035 0.795 2.915 0.795 2.915 0.635 2.515 0.635 2.515 0.415 2.195 0.415 2.195 0.685 2.255 0.685 2.255 0.745 2.135 0.745 2.135 0.355 2.575 0.355 2.575 0.575 2.915 0.575 2.915 0.355 3.745 0.355 ;
      POLYGON 3.195 1.305 3.135 1.305 3.135 0.955 2.515 0.955 2.515 0.895 3.135 0.895 3.135 0.575 3.075 0.575 3.075 0.515 3.195 0.515 ;
      POLYGON 3.085 1.465 2.965 1.465 2.965 1.305 1.685 1.305 1.685 1.15 0.84 1.15 0.84 0.57 0.96 0.57 0.96 0.63 0.9 0.63 0.9 1.09 1.685 1.09 1.685 0.825 1.625 0.825 1.625 0.765 1.745 0.765 1.745 1.245 2.005 1.245 2.005 0.855 2.065 0.855 2.065 1.245 3.025 1.245 3.025 1.405 3.085 1.405 ;
      POLYGON 2.815 0.795 2.415 0.795 2.415 1.115 2.295 1.115 2.295 1.055 2.355 1.055 2.355 0.575 2.295 0.575 2.295 0.515 2.415 0.515 2.415 0.735 2.815 0.735 ;
      POLYGON 1.905 1.145 1.845 1.145 1.845 0.665 1.365 0.665 1.365 0.83 1.305 0.83 1.305 0.605 1.845 0.605 1.845 0.485 1.905 0.485 ;
      POLYGON 1.525 0.99 1.085 0.99 1.085 0.93 1.145 0.93 1.145 0.47 0.735 0.47 0.735 0.65 0.56 0.65 0.56 0.79 0.44 0.79 0.44 0.59 0.675 0.59 0.675 0.41 1.205 0.41 1.205 0.93 1.465 0.93 1.465 0.855 1.525 0.855 ;
  END
END SMDFFHQX2

MACRO SMDFFHQX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SMDFFHQX4 0 0 ;
  SIZE 6.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.019802 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.39 0.765 6.33 0.765 6.33 0.705 5.66 0.705 5.66 0.99 5.6 0.99 5.6 0.645 6.235 0.645 6.235 0.625 6.365 0.625 6.365 0.645 6.39 0.645 ;
    END
  END S0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.23 0.885 6.165 0.885 6.165 1.085 5.93 1.085 5.93 0.805 6.23 0.805 ;
    END
  END D1
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.26 0.455 5.34 0.955 ;
    END
  END D0
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.82838275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.06 0.455 5.14 0.955 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.105 0.92 3.86 0.92 3.86 0.79 4.025 0.79 4.025 0.585 4.105 0.585 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.42 0.34 0.92 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5408 LAYER Metal1 ;
    ANTENNADIFFAREA 4.5142 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.400275 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.8459185 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 68.7877085 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.13 1.05 0.46 1.05 0.46 0.79 0.53 0.79 0.53 0.535 0.59 0.535 0.59 0.99 0.895 0.99 0.895 0.65 0.94 0.65 0.94 0.535 1 0.535 1 0.71 0.955 0.71 0.955 0.99 1.13 0.99 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.8 1.77 0 1.77 0 1.65 0.335 1.65 0.335 1.51 0.395 1.51 0.395 1.65 0.775 1.65 0.775 1.34 0.895 1.34 0.895 1.4 0.835 1.4 0.835 1.65 1.245 1.65 1.245 1.34 1.365 1.34 1.365 1.4 1.305 1.4 1.305 1.65 1.715 1.65 1.715 1.34 1.835 1.34 1.835 1.4 1.775 1.4 1.775 1.65 2.835 1.65 2.835 1.34 2.955 1.34 2.955 1.4 2.895 1.4 2.895 1.65 4.015 1.65 4.015 1.24 4.075 1.24 4.075 1.65 5.25 1.65 5.25 1.215 5.31 1.215 5.31 1.65 6.015 1.65 6.015 1.36 6.075 1.36 6.075 1.65 6.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.8 0.06 6.18 0.06 6.18 0.47 6.12 0.47 6.12 0.06 5.3 0.06 5.3 0.355 5.24 0.355 5.24 0.06 4.145 0.06 4.145 0.485 4.085 0.485 4.085 0.06 2.955 0.06 2.955 0.17 2.835 0.17 2.835 0.06 1.615 0.06 1.615 0.34 1.675 0.34 1.675 0.4 1.555 0.4 1.555 0.06 1.205 0.06 1.205 0.515 1.145 0.515 1.145 0.06 0.795 0.06 0.795 0.515 0.735 0.515 0.735 0.06 0.355 0.06 0.355 0.2 0.295 0.2 0.295 0.06 0 0.06 0 -0.06 6.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 6.55 0.925 6.465 0.925 6.465 1.305 6.405 1.305 6.405 1.245 5.77 1.245 5.77 0.93 5.83 0.93 5.83 1.185 6.405 1.185 6.405 0.865 6.49 0.865 6.49 0.375 6.55 0.375 ;
      POLYGON 5.87 0.495 5.5 0.495 5.5 1.09 5.67 1.09 5.67 1.48 5.61 1.48 5.61 1.15 5.44 1.15 5.44 1.115 4.745 1.115 4.745 1.175 4.685 1.175 4.685 1.055 4.79 1.055 4.79 0.5 4.85 0.5 4.85 1.055 5.44 1.055 5.44 0.435 5.81 0.435 5.81 0.375 5.87 0.375 ;
      POLYGON 5.105 1.335 4.525 1.335 4.525 0.86 4.425 0.86 4.425 0.92 4.365 0.92 4.365 0.8 4.63 0.8 4.63 0.235 5.075 0.235 5.075 0.355 5.015 0.355 5.015 0.295 4.69 0.295 4.69 0.86 4.585 0.86 4.585 1.275 4.985 1.275 4.985 1.215 5.105 1.215 ;
      POLYGON 4.53 0.7 4.265 0.7 4.265 1.02 4.425 1.02 4.425 1.36 4.365 1.36 4.365 1.08 3.65 1.08 3.65 0.51 3.77 0.51 3.77 0.57 3.71 0.57 3.71 1.02 4.205 1.02 4.205 0.64 4.47 0.64 4.47 0.5 4.53 0.5 ;
      POLYGON 3.94 0.485 3.88 0.485 3.88 0.4 3.55 0.4 3.55 1.19 3.9 1.19 3.9 1.25 3.49 1.25 3.49 0.4 3.17 0.4 3.17 0.66 3.19 0.66 3.19 0.78 3.11 0.78 3.11 0.41 2.355 0.41 2.355 0.67 2.47 0.67 2.47 0.73 2.295 0.73 2.295 0.35 3.11 0.35 3.11 0.34 3.94 0.34 ;
      POLYGON 3.39 1.24 3.33 1.24 3.33 0.94 2.79 0.94 2.79 0.88 2.73 0.88 2.73 0.82 2.85 0.82 2.85 0.88 3.33 0.88 3.33 0.56 3.27 0.56 3.27 0.5 3.39 0.5 ;
      POLYGON 3.28 1.4 3.16 1.4 3.16 1.24 2.37 1.24 2.37 1.27 1.99 1.27 1.99 1.24 0.1 1.24 0.1 0.535 0.16 0.535 0.16 1.18 1.85 1.18 1.85 0.66 1.91 0.66 1.91 1.18 2.05 1.18 2.05 1.21 2.31 1.21 2.31 0.89 2.17 0.89 2.17 0.83 2.37 0.83 2.37 1.18 3.22 1.18 3.22 1.34 3.28 1.34 ;
      POLYGON 3.01 0.77 2.95 0.77 2.95 0.71 2.63 0.71 2.63 1.08 2.57 1.08 2.57 0.57 2.455 0.57 2.455 0.51 2.63 0.51 2.63 0.65 3.01 0.65 ;
      POLYGON 2.21 1.11 2.15 1.11 2.15 1.05 2.01 1.05 2.01 0.56 1.57 0.56 1.57 0.76 1.51 0.76 1.51 0.5 2.01 0.5 2.01 0.44 2.07 0.44 2.07 0.99 2.21 0.99 ;
      POLYGON 1.75 0.92 1.41 0.92 1.41 1.02 1.6 1.02 1.6 1.08 1.35 1.08 1.35 0.865 1.055 0.865 1.055 0.805 1.35 0.805 1.35 0.48 1.41 0.48 1.41 0.86 1.69 0.86 1.69 0.66 1.75 0.66 ;
  END
END SMDFFHQX4

MACRO SMDFFHQX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SMDFFHQX8 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN S0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.54785475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.715 0.765 7.655 0.765 7.655 0.705 7.08 0.705 7.08 0.755 6.92 0.755 6.92 0.945 6.8 0.945 6.8 0.885 6.86 0.885 6.86 0.695 7.02 0.695 7.02 0.645 7.035 0.645 7.035 0.625 7.205 0.625 7.205 0.645 7.715 0.645 ;
    END
  END S0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.555 0.885 7.375 0.885 7.375 1.01 7.18 1.01 7.18 0.805 7.555 0.805 ;
    END
  END D1
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.54 0.995 6.42 0.995 6.42 0.885 6.46 0.885 6.46 0.535 6.54 0.535 ;
    END
  END D0
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.82838275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.34 0.73 6.32 0.73 6.32 1.005 6.24 1.005 6.24 0.65 6.26 0.65 6.26 0.525 6.34 0.525 ;
    END
  END SE
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.02925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.948718 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.395 1.01 5.26 1.01 5.26 0.565 5.34 0.565 5.34 0.86 5.395 0.86 ;
    END
  END SI
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.93 0.895 2.605 0.895 2.605 0.815 2.82 0.815 2.82 0.64 2.93 0.64 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.39425 LAYER Metal1 ;
    ANTENNADIFFAREA 5.394675 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.557775 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.87817675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 62.2509075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.37 0.65 1.325 0.65 1.325 0.9 1.37 0.9 1.37 1.345 1.31 1.345 1.31 0.96 1.265 0.96 1.265 0.8 0.96 0.8 0.96 1.345 0.9 1.345 0.9 0.66 0.55 0.66 0.55 1.345 0.49 1.345 0.49 0.66 0.14 0.66 0.14 1.345 0.08 1.345 0.08 0.73 0.06 0.73 0.06 0.6 0.08 0.6 0.08 0.54 0.14 0.54 0.14 0.6 0.49 0.6 0.49 0.54 0.55 0.54 0.55 0.6 0.9 0.6 0.9 0.54 0.96 0.54 0.96 0.74 1.265 0.74 1.265 0.59 1.31 0.59 1.31 0.53 1.37 0.53 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 1.77 0 1.77 0 1.65 0.285 1.65 0.285 0.9 0.345 0.9 0.345 1.65 0.695 1.65 0.695 0.9 0.755 0.9 0.755 1.65 1.105 1.65 1.105 0.9 1.165 0.9 1.165 1.65 1.515 1.65 1.515 0.955 1.575 0.955 1.575 1.65 1.925 1.65 1.925 1.055 1.985 1.055 1.985 1.65 2.98 1.65 2.98 1.315 3.04 1.315 3.04 1.65 4.12 1.65 4.12 1.365 4.24 1.365 4.24 1.425 4.18 1.425 4.18 1.65 5.42 1.65 5.42 1.27 5.48 1.27 5.48 1.65 6.55 1.65 6.55 1.285 6.61 1.285 6.61 1.65 7.36 1.65 7.36 1.285 7.42 1.285 7.42 1.65 8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 0.06 7.42 0.06 7.42 0.545 7.36 0.545 7.36 0.06 6.625 0.06 6.625 0.435 6.565 0.435 6.565 0.06 5.48 0.06 5.48 0.465 5.42 0.465 5.42 0.06 4.29 0.06 4.29 0.365 4.17 0.365 4.17 0.305 4.23 0.305 4.23 0.06 3.015 0.06 3.015 0.22 2.895 0.22 2.895 0.16 2.955 0.16 2.955 0.06 1.985 0.06 1.985 0.485 1.925 0.485 1.925 0.06 1.575 0.06 1.575 0.485 1.515 0.485 1.515 0.06 1.165 0.06 1.165 0.485 1.105 0.485 1.105 0.06 0.755 0.06 0.755 0.485 0.695 0.485 0.695 0.06 0.345 0.06 0.345 0.485 0.285 0.485 0.285 0.06 0 0.06 0 -0.06 8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.875 1.17 7.79 1.17 7.79 1.23 7.73 1.23 7.73 1.17 7.02 1.17 7.02 0.855 7.08 0.855 7.08 1.11 7.815 1.11 7.815 0.45 7.875 0.45 ;
      POLYGON 7.11 0.525 6.92 0.525 6.92 0.595 6.7 0.595 6.7 1.105 6.92 1.105 6.92 1.405 6.86 1.405 6.86 1.165 6.05 1.165 6.05 1 6.08 1 6.08 0.375 6.2 0.375 6.2 0.435 6.14 0.435 6.14 1.105 6.64 1.105 6.64 0.535 6.86 0.535 6.86 0.465 7.05 0.465 7.05 0.405 7.11 0.405 ;
      POLYGON 6.42 0.425 6.3 0.425 6.3 0.275 5.98 0.275 5.98 0.89 5.95 0.89 5.95 1.265 6.405 1.265 6.405 1.385 6.345 1.385 6.345 1.325 5.89 1.325 5.89 0.89 5.715 0.89 5.715 0.95 5.655 0.95 5.655 0.83 5.92 0.83 5.92 0.215 6.36 0.215 6.36 0.365 6.42 0.365 ;
      POLYGON 5.82 0.575 5.64 0.575 5.64 0.625 5.555 0.625 5.555 1.11 5.79 1.11 5.79 1.39 5.73 1.39 5.73 1.17 5.045 1.17 5.045 1.23 4.985 1.23 4.985 0.505 5.105 0.505 5.105 0.565 5.045 0.565 5.045 1.11 5.495 1.11 5.495 0.565 5.58 0.565 5.58 0.515 5.82 0.515 ;
      POLYGON 5.305 1.36 5.205 1.36 5.205 1.39 4.825 1.39 4.825 0.405 4.505 0.405 4.505 0.665 4.565 0.665 4.565 0.725 4.445 0.725 4.445 0.525 4.01 0.525 4.01 0.345 3.69 0.345 3.69 0.605 3.75 0.605 3.75 0.77 3.69 0.77 3.69 0.665 3.63 0.665 3.63 0.285 4.07 0.285 4.07 0.465 4.445 0.465 4.445 0.345 5.275 0.345 5.275 0.465 5.215 0.465 5.215 0.405 4.885 0.405 4.885 1.33 5.145 1.33 5.145 1.3 5.305 1.3 ;
      POLYGON 4.725 1.235 4.665 1.235 4.665 0.885 4.075 0.885 4.075 0.845 4.015 0.845 4.015 0.785 4.135 0.785 4.135 0.825 4.665 0.825 4.665 0.565 4.605 0.565 4.605 0.505 4.725 0.505 ;
      POLYGON 4.565 1.395 4.505 1.395 4.505 1.265 3.2 1.265 3.2 0.54 2.505 0.54 2.505 0.995 2.835 0.995 2.835 1.055 2.445 1.055 2.445 0.48 3.26 0.48 3.26 1.205 3.535 1.205 3.535 0.885 3.52 0.885 3.52 0.765 3.58 0.765 3.58 0.825 3.595 0.825 3.595 1.205 4.565 1.205 ;
      POLYGON 4.345 0.725 4.225 0.725 4.225 0.685 3.91 0.685 3.91 1.045 3.85 1.045 3.85 0.505 3.79 0.505 3.79 0.445 3.91 0.445 3.91 0.625 4.285 0.625 4.285 0.665 4.345 0.665 ;
      POLYGON 3.435 1.105 3.375 1.105 3.375 1.045 3.36 1.045 3.36 0.38 2.145 0.38 2.145 0.795 2.085 0.795 2.085 0.32 3.42 0.32 3.42 0.985 3.435 0.985 ;
      POLYGON 3.09 1.215 2.19 1.215 2.19 1.345 2.13 1.345 2.13 1.055 2.245 1.055 2.245 0.955 1.78 0.955 1.78 1.345 1.72 1.345 1.72 0.805 1.425 0.805 1.425 0.745 1.72 0.745 1.72 0.505 1.78 0.505 1.78 0.895 2.245 0.895 2.245 0.505 2.305 0.505 2.305 1.155 3.03 1.155 3.03 0.73 3.09 0.73 ;
  END
END SMDFFHQX8

MACRO SPDFF2RX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SPDFF2RX1 0 0 ;
  SIZE 10.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1511 LAYER Metal1 ;
    ANTENNADIFFAREA 10.171375 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4572 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.4538495 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 99.816273 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.14 0.96 10.09 0.96 10.09 1.11 9.96 1.11 9.96 1.05 9.995 1.05 9.995 0.54 10.07 0.54 10.07 0.6 10.075 0.6 10.075 0.76 10.14 0.76 ;
    END
  END Q2
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1511 LAYER Metal1 ;
    ANTENNADIFFAREA 10.233375 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4572 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.4538495 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 99.816273 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.74 1.11 10.61 1.11 10.61 1.05 10.645 1.05 10.645 0.54 10.74 0.54 ;
    END
  END Q2N
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.14 0.875 7.06 0.875 7.06 0.775 7.015 0.775 7.015 0.62 7.14 0.62 ;
    END
  END D2
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7513 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0648 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.59413575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 108.47222225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.735 1.35 7.735 1.35 7.735 1.375 7.335 1.375 7.335 1.35 5.75 1.35 5.75 1.465 5.46 1.465 5.46 1.35 3.465 1.35 3.465 1.375 3.065 1.375 3.065 1.35 0.065 1.35 0.065 1.29 3.125 1.29 3.125 1.315 3.41 1.315 3.41 1.29 7.39 1.29 7.39 1.315 7.675 1.315 7.675 1.29 10.735 1.29 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0648 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 60.83333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.735 0.41 6.57 0.41 6.57 0.7 6.835 0.7 6.835 0.865 6.775 0.865 6.775 0.76 6.51 0.76 6.51 0.41 6.145 0.41 6.145 0.895 6.06 0.895 6.06 0.41 4.74 0.41 4.74 0.895 4.655 0.895 4.655 0.41 4.29 0.41 4.29 0.76 4.025 0.76 4.025 0.865 3.965 0.865 3.965 0.7 4.23 0.7 4.23 0.41 0.065 0.41 0.065 0.35 10.735 0.35 ;
    END
  END SE
  PIN SI2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.235 0.625 6.41 0.77 ;
    END
  END SI2
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1511 LAYER Metal1 ;
    ANTENNADIFFAREA 8.651875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4572 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.4538495 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 99.816273 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.84 1.11 0.71 1.11 0.71 0.96 0.66 0.96 0.66 0.76 0.725 0.76 0.725 0.6 0.73 0.6 0.73 0.54 0.805 0.54 0.805 1.05 0.84 1.05 ;
    END
  END Q1
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.1511 LAYER Metal1 ;
    ANTENNADIFFAREA 8.603325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4572 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.4538495 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 99.816273 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.19 1.11 0.06 1.11 0.06 0.54 0.155 0.54 0.155 1.05 0.19 1.05 ;
    END
  END Q1N
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.785 0.775 3.74 0.775 3.74 0.875 3.66 0.875 3.66 0.62 3.785 0.62 ;
    END
  END D1
  PIN SI1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.39 0.625 4.565 0.77 ;
    END
  END SI1
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.445 0.77 5.625 0.92 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.8 1.77 0 1.77 0 1.65 0.3 1.65 0.3 1.54 0.42 1.54 0.42 1.65 0.955 1.65 0.955 1.54 1.075 1.54 1.075 1.65 1.53 1.65 1.53 1.54 1.65 1.54 1.65 1.65 2.445 1.65 2.445 1.54 2.565 1.54 2.565 1.65 2.795 1.65 2.795 1.54 2.915 1.54 2.915 1.65 3.675 1.65 3.675 1.54 3.795 1.54 3.795 1.65 4.465 1.65 4.465 1.54 4.585 1.54 4.585 1.65 5.33 1.65 5.33 1.54 5.45 1.54 5.45 1.65 6.215 1.65 6.215 1.54 6.335 1.54 6.335 1.65 7.005 1.65 7.005 1.54 7.125 1.54 7.125 1.65 7.885 1.65 7.885 1.54 8.005 1.54 8.005 1.65 8.235 1.65 8.235 1.54 8.355 1.54 8.355 1.65 9.15 1.65 9.15 1.54 9.27 1.54 9.27 1.65 9.725 1.65 9.725 1.54 9.845 1.54 9.845 1.65 10.38 1.65 10.38 1.54 10.5 1.54 10.5 1.65 10.8 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.8 0.06 10.5 0.06 10.5 0.17 10.38 0.17 10.38 0.06 9.895 0.06 9.895 0.17 9.775 0.17 9.775 0.06 9.27 0.06 9.27 0.17 9.15 0.17 9.15 0.06 8.255 0.06 8.255 0.17 8.135 0.17 8.135 0.06 7.15 0.06 7.15 0.17 7.03 0.17 7.03 0.06 6.335 0.06 6.335 0.17 6.215 0.17 6.215 0.06 5.45 0.06 5.45 0.17 5.325 0.17 5.325 0.06 4.585 0.06 4.585 0.17 4.465 0.17 4.465 0.06 3.77 0.06 3.77 0.17 3.65 0.17 3.65 0.06 2.665 0.06 2.665 0.17 2.545 0.17 2.545 0.06 1.65 0.06 1.65 0.17 1.53 0.17 1.53 0.06 1.025 0.06 1.025 0.17 0.905 0.17 0.905 0.06 0.42 0.06 0.42 0.17 0.3 0.17 0.3 0.06 0 0.06 0 -0.06 10.8 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 10.735 0.29 0.065 0.29 0.065 0.23 4.66 0.23 4.66 0.205 4.8 0.205 4.8 0.23 6 0.23 6 0.205 6.14 0.205 6.14 0.23 10.735 0.23 ;
      POLYGON 10.735 1.23 7.615 1.23 7.615 1.255 7.45 1.255 7.45 1.23 3.35 1.23 3.35 1.255 3.185 1.255 3.185 1.23 0.065 1.23 0.065 1.17 1.835 1.17 1.835 0.665 1.895 0.665 1.895 1.17 2.165 1.17 2.165 0.865 2.105 0.865 2.105 0.805 2.225 0.805 2.225 1.17 4.64 1.17 4.64 1.15 4.78 1.15 4.78 1.17 5.3 1.17 5.3 0.895 5.26 0.895 5.26 0.495 5.36 0.495 5.36 0.625 5.565 0.625 5.565 0.505 5.625 0.505 5.625 0.705 5.36 0.705 5.36 1.005 5.655 1.005 5.655 1.065 5.36 1.065 5.36 1.17 6.02 1.17 6.02 1.15 6.16 1.15 6.16 1.17 8.575 1.17 8.575 0.805 8.695 0.805 8.695 0.865 8.635 0.865 8.635 1.17 8.905 1.17 8.905 0.665 8.965 0.665 8.965 1.17 10.735 1.17 ;
      POLYGON 10.73 1.48 7.84 1.48 7.84 1.495 7.22 1.495 7.22 1.48 7.005 1.48 7.005 1.42 7.275 1.42 7.275 1.435 7.78 1.435 7.78 1.42 10.73 1.42 ;
      POLYGON 10.545 0.84 10.29 0.84 10.29 1.02 10.21 1.02 10.21 0.54 10.29 0.54 10.29 0.76 10.545 0.76 ;
      POLYGON 9.925 0.82 9.645 0.82 9.645 1.1 9.075 1.1 9.075 0.68 9.135 0.68 9.135 1.04 9.585 1.04 9.585 0.485 9.645 0.485 9.645 0.76 9.925 0.76 ;
      POLYGON 9.515 0.825 9.455 0.825 9.455 0.66 9.4 0.66 9.4 0.575 8.82 0.575 8.82 1.055 8.76 1.055 8.76 0.575 8.71 0.575 8.71 0.495 9.46 0.495 9.46 0.6 9.515 0.6 ;
      RECT 9.235 0.735 9.395 0.96 ;
      POLYGON 8.54 0.575 8.51 0.575 8.51 1.055 8.45 1.055 8.45 0.74 7.855 0.74 7.855 0.68 8.45 0.68 8.45 0.575 8.42 0.575 8.42 0.515 8.54 0.515 ;
      POLYGON 8.37 0.86 7.52 0.86 7.52 1.045 7.46 1.045 7.46 0.8 7.645 0.8 7.645 0.575 7.61 0.575 7.61 0.515 7.74 0.515 7.74 0.575 7.705 0.575 7.705 0.8 8.37 0.8 ;
      RECT 7.635 0.95 8.135 1.03 ;
      POLYGON 7.53 0.575 7.5 0.575 7.5 0.73 7.4 0.73 7.4 0.95 7.315 0.95 7.315 1.065 6.615 1.065 6.615 1.005 6.895 1.005 6.895 0.54 6.655 0.54 6.655 0.48 6.955 0.48 6.955 1.005 7.255 1.005 7.255 0.89 7.34 0.89 7.34 0.67 7.44 0.67 7.44 0.575 7.41 0.575 7.41 0.515 7.53 0.515 ;
      POLYGON 6.67 0.905 6.315 0.905 6.315 1.065 5.925 1.065 5.925 0.51 5.985 0.51 5.985 1.005 6.255 1.005 6.255 0.845 6.67 0.845 ;
      RECT 5.925 1.42 6.495 1.48 ;
      POLYGON 5.2 1.1 5.06 1.1 5.06 0.77 5.14 0.77 5.14 0.495 5.2 0.495 ;
      POLYGON 4.875 1.065 4.485 1.065 4.485 0.905 4.13 0.905 4.13 0.845 4.545 0.845 4.545 1.005 4.815 1.005 4.815 0.51 4.875 0.51 ;
      RECT 4.305 1.42 4.875 1.48 ;
      POLYGON 4.185 1.065 3.485 1.065 3.485 0.95 3.4 0.95 3.4 0.73 3.3 0.73 3.3 0.575 3.27 0.575 3.27 0.515 3.39 0.515 3.39 0.575 3.36 0.575 3.36 0.67 3.46 0.67 3.46 0.89 3.545 0.89 3.545 1.005 3.845 1.005 3.845 0.48 4.145 0.48 4.145 0.54 3.905 0.54 3.905 1.005 4.185 1.005 ;
      POLYGON 3.795 1.48 3.58 1.48 3.58 1.495 2.96 1.495 2.96 1.48 0.07 1.48 0.07 1.42 3.02 1.42 3.02 1.435 3.525 1.435 3.525 1.42 3.795 1.42 ;
      POLYGON 3.34 1.045 3.28 1.045 3.28 0.86 2.43 0.86 2.43 0.8 3.095 0.8 3.095 0.575 3.06 0.575 3.06 0.515 3.19 0.515 3.19 0.575 3.155 0.575 3.155 0.8 3.34 0.8 ;
      RECT 2.665 0.95 3.165 1.03 ;
      POLYGON 2.945 0.74 2.35 0.74 2.35 1.055 2.29 1.055 2.29 0.575 2.26 0.575 2.26 0.515 2.38 0.515 2.38 0.575 2.35 0.575 2.35 0.68 2.945 0.68 ;
      POLYGON 2.09 0.575 2.04 0.575 2.04 1.055 1.98 1.055 1.98 0.575 1.4 0.575 1.4 0.66 1.345 0.66 1.345 0.825 1.285 0.825 1.285 0.6 1.34 0.6 1.34 0.495 2.09 0.495 ;
      POLYGON 1.725 1.1 1.155 1.1 1.155 0.82 0.875 0.82 0.875 0.76 1.155 0.76 1.155 0.485 1.215 0.485 1.215 1.04 1.665 1.04 1.665 0.68 1.725 0.68 ;
      RECT 1.405 0.735 1.565 0.96 ;
      POLYGON 0.59 1.02 0.51 1.02 0.51 0.84 0.255 0.84 0.255 0.76 0.51 0.76 0.51 0.54 0.59 0.54 ;
  END
END SPDFF2RX1

MACRO SPDFF2RX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SPDFF2RX2 0 0 ;
  SIZE 12 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3917 LAYER Metal1 ;
    ANTENNADIFFAREA 11.986325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.58815 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.86746575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 76.67431775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.585 0.54 10.74 1.11 ;
    END
  END Q2
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.74 0.875 7.66 0.875 7.66 0.775 7.615 0.775 7.615 0.62 7.74 0.62 ;
    END
  END D2
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3917 LAYER Metal1 ;
    ANTENNADIFFAREA 11.673125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.58815 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.86746575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 76.67431775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.455 0.54 11.595 1.11 ;
    END
  END Q2N
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.6247 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.07875 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.9326985 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 73.1809525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.28 1.35 8.335 1.35 8.335 1.375 7.935 1.375 7.935 1.35 6.35 1.35 6.35 1.465 6.06 1.465 6.06 1.35 4.065 1.35 4.065 1.375 3.665 1.375 3.665 1.35 1.72 1.35 1.72 1.29 3.725 1.29 3.725 1.315 4.01 1.315 4.01 1.29 7.99 1.29 7.99 1.315 8.275 1.315 8.275 1.29 10.28 1.29 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0648 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 51.06481475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 10.28 0.41 7.17 0.41 7.17 0.7 7.435 0.7 7.435 0.865 7.375 0.865 7.375 0.76 7.11 0.76 7.11 0.41 6.745 0.41 6.745 0.895 6.66 0.895 6.66 0.41 5.34 0.41 5.34 0.895 5.255 0.895 5.255 0.41 4.89 0.41 4.89 0.76 4.625 0.76 4.625 0.865 4.565 0.865 4.565 0.7 4.83 0.7 4.83 0.41 1.72 0.41 1.72 0.35 10.28 0.35 ;
    END
  END SE
  PIN SI2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.835 0.625 7.01 0.77 ;
    END
  END SI2
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3917 LAYER Metal1 ;
    ANTENNADIFFAREA 9.920025 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.58815 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.86746575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 76.67431775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.54 1.415 1.11 ;
    END
  END Q1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.385 0.775 4.34 0.775 4.34 0.875 4.26 0.875 4.26 0.62 4.385 0.62 ;
    END
  END D1
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.3917 LAYER Metal1 ;
    ANTENNADIFFAREA 9.896075 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.58815 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.86746575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 76.67431775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.405 0.54 0.545 1.11 ;
    END
  END Q1N
  PIN SI1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.99 0.625 5.165 0.77 ;
    END
  END SI1
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.045 0.77 6.225 0.92 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 12 1.77 0 1.77 0 1.65 0.24 1.65 0.24 1.54 0.36 1.54 0.36 1.65 0.61 1.65 0.61 1.54 0.765 1.54 0.765 1.65 1.065 1.65 1.065 1.54 1.185 1.54 1.185 1.65 1.555 1.65 1.555 1.54 1.675 1.54 1.675 1.65 2.13 1.65 2.13 1.54 2.25 1.54 2.25 1.65 3.045 1.65 3.045 1.54 3.165 1.54 3.165 1.65 3.395 1.65 3.395 1.54 3.515 1.54 3.515 1.65 4.275 1.65 4.275 1.54 4.395 1.54 4.395 1.65 5.065 1.65 5.065 1.54 5.185 1.54 5.185 1.65 5.93 1.65 5.93 1.54 6.05 1.54 6.05 1.65 6.815 1.65 6.815 1.54 6.935 1.54 6.935 1.65 7.605 1.65 7.605 1.54 7.725 1.54 7.725 1.65 8.485 1.65 8.485 1.54 8.605 1.54 8.605 1.65 8.835 1.65 8.835 1.54 8.955 1.54 8.955 1.65 9.75 1.65 9.75 1.54 9.87 1.54 9.87 1.65 10.325 1.65 10.325 1.54 10.445 1.54 10.445 1.65 10.815 1.65 10.815 1.54 10.935 1.54 10.935 1.65 11.235 1.65 11.235 1.54 11.39 1.54 11.39 1.65 11.64 1.65 11.64 1.54 11.76 1.54 11.76 1.65 12 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 12 0.06 11.76 0.06 11.76 0.17 11.64 0.17 11.64 0.06 11.39 0.06 11.39 0.17 11.27 0.17 11.27 0.06 10.935 0.06 10.935 0.17 10.815 0.17 10.815 0.06 10.495 0.06 10.495 0.17 10.375 0.17 10.375 0.06 9.87 0.06 9.87 0.17 9.75 0.17 9.75 0.06 8.855 0.06 8.855 0.17 8.735 0.17 8.735 0.06 7.75 0.06 7.75 0.17 7.63 0.17 7.63 0.06 6.935 0.06 6.935 0.17 6.815 0.17 6.815 0.06 6.05 0.06 6.05 0.17 5.925 0.17 5.925 0.06 5.185 0.06 5.185 0.17 5.065 0.17 5.065 0.06 4.37 0.06 4.37 0.17 4.25 0.17 4.25 0.06 3.265 0.06 3.265 0.17 3.145 0.17 3.145 0.06 2.25 0.06 2.25 0.17 2.13 0.17 2.13 0.06 1.625 0.06 1.625 0.17 1.505 0.17 1.505 0.06 1.185 0.06 1.185 0.17 1.065 0.17 1.065 0.06 0.73 0.06 0.73 0.17 0.61 0.17 0.61 0.06 0.36 0.06 0.36 0.17 0.24 0.17 0.24 0.06 0 0.06 0 -0.06 12 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 11.37 0.85 11.31 0.85 11.31 0.82 11.145 0.82 11.145 1.02 11.065 1.02 11.065 0.54 11.145 0.54 11.145 0.76 11.31 0.76 11.31 0.725 11.37 0.725 ;
      POLYGON 10.525 0.82 10.245 0.82 10.245 1.1 9.675 1.1 9.675 0.68 9.735 0.68 9.735 1.04 10.185 1.04 10.185 0.485 10.245 0.485 10.245 0.76 10.525 0.76 ;
      POLYGON 10.28 0.29 1.72 0.29 1.72 0.23 5.26 0.23 5.26 0.205 5.4 0.205 5.4 0.23 6.6 0.23 6.6 0.205 6.74 0.205 6.74 0.23 10.28 0.23 ;
      POLYGON 10.28 1.23 8.215 1.23 8.215 1.255 8.05 1.255 8.05 1.23 3.95 1.23 3.95 1.255 3.785 1.255 3.785 1.23 1.72 1.23 1.72 1.17 2.435 1.17 2.435 0.665 2.495 0.665 2.495 1.17 2.765 1.17 2.765 0.865 2.705 0.865 2.705 0.805 2.825 0.805 2.825 1.17 5.24 1.17 5.24 1.15 5.38 1.15 5.38 1.17 5.9 1.17 5.9 0.895 5.86 0.895 5.86 0.495 5.96 0.495 5.96 0.625 6.165 0.625 6.165 0.505 6.225 0.505 6.225 0.705 5.96 0.705 5.96 1.005 6.255 1.005 6.255 1.065 5.96 1.065 5.96 1.17 6.62 1.17 6.62 1.15 6.76 1.15 6.76 1.17 9.175 1.17 9.175 0.805 9.295 0.805 9.295 0.865 9.235 0.865 9.235 1.17 9.505 1.17 9.505 0.665 9.565 0.665 9.565 1.17 10.28 1.17 ;
      POLYGON 10.275 1.48 8.44 1.48 8.44 1.495 7.82 1.495 7.82 1.48 7.605 1.48 7.605 1.42 7.875 1.42 7.875 1.435 8.38 1.435 8.38 1.42 10.275 1.42 ;
      POLYGON 10.115 0.825 10.055 0.825 10.055 0.66 10 0.66 10 0.575 9.42 0.575 9.42 1.055 9.36 1.055 9.36 0.575 9.31 0.575 9.31 0.495 10.06 0.495 10.06 0.6 10.115 0.6 ;
      RECT 9.835 0.735 9.995 0.96 ;
      POLYGON 9.14 0.575 9.11 0.575 9.11 1.055 9.05 1.055 9.05 0.74 8.455 0.74 8.455 0.68 9.05 0.68 9.05 0.575 9.02 0.575 9.02 0.515 9.14 0.515 ;
      POLYGON 8.97 0.86 8.12 0.86 8.12 1.045 8.06 1.045 8.06 0.8 8.245 0.8 8.245 0.575 8.21 0.575 8.21 0.515 8.34 0.515 8.34 0.575 8.305 0.575 8.305 0.8 8.97 0.8 ;
      RECT 8.235 0.95 8.735 1.03 ;
      POLYGON 8.13 0.575 8.1 0.575 8.1 0.73 8 0.73 8 0.95 7.915 0.95 7.915 1.065 7.215 1.065 7.215 1.005 7.495 1.005 7.495 0.54 7.255 0.54 7.255 0.48 7.555 0.48 7.555 1.005 7.855 1.005 7.855 0.89 7.94 0.89 7.94 0.67 8.04 0.67 8.04 0.575 8.01 0.575 8.01 0.515 8.13 0.515 ;
      POLYGON 7.27 0.905 6.915 0.905 6.915 1.065 6.525 1.065 6.525 0.51 6.585 0.51 6.585 1.005 6.855 1.005 6.855 0.845 7.27 0.845 ;
      RECT 6.525 1.42 7.095 1.48 ;
      POLYGON 5.8 1.1 5.66 1.1 5.66 0.77 5.74 0.77 5.74 0.495 5.8 0.495 ;
      POLYGON 5.475 1.065 5.085 1.065 5.085 0.905 4.73 0.905 4.73 0.845 5.145 0.845 5.145 1.005 5.415 1.005 5.415 0.51 5.475 0.51 ;
      RECT 4.905 1.42 5.475 1.48 ;
      POLYGON 4.785 1.065 4.085 1.065 4.085 0.95 4 0.95 4 0.73 3.9 0.73 3.9 0.575 3.87 0.575 3.87 0.515 3.99 0.515 3.99 0.575 3.96 0.575 3.96 0.67 4.06 0.67 4.06 0.89 4.145 0.89 4.145 1.005 4.445 1.005 4.445 0.48 4.745 0.48 4.745 0.54 4.505 0.54 4.505 1.005 4.785 1.005 ;
      POLYGON 4.395 1.48 4.18 1.48 4.18 1.495 3.56 1.495 3.56 1.48 1.725 1.48 1.725 1.42 3.62 1.42 3.62 1.435 4.125 1.435 4.125 1.42 4.395 1.42 ;
      POLYGON 3.94 1.045 3.88 1.045 3.88 0.86 3.03 0.86 3.03 0.8 3.695 0.8 3.695 0.575 3.66 0.575 3.66 0.515 3.79 0.515 3.79 0.575 3.755 0.575 3.755 0.8 3.94 0.8 ;
      RECT 3.265 0.95 3.765 1.03 ;
      POLYGON 3.545 0.74 2.95 0.74 2.95 1.055 2.89 1.055 2.89 0.575 2.86 0.575 2.86 0.515 2.98 0.515 2.98 0.575 2.95 0.575 2.95 0.68 3.545 0.68 ;
      POLYGON 2.69 0.575 2.64 0.575 2.64 1.055 2.58 1.055 2.58 0.575 2 0.575 2 0.66 1.945 0.66 1.945 0.825 1.885 0.825 1.885 0.6 1.94 0.6 1.94 0.495 2.69 0.495 ;
      POLYGON 2.325 1.1 1.755 1.1 1.755 0.82 1.475 0.82 1.475 0.76 1.755 0.76 1.755 0.485 1.815 0.485 1.815 1.04 2.265 1.04 2.265 0.68 2.325 0.68 ;
      RECT 2.005 0.735 2.165 0.96 ;
      POLYGON 0.935 1.02 0.855 1.02 0.855 0.82 0.69 0.82 0.69 0.85 0.63 0.85 0.63 0.725 0.69 0.725 0.69 0.76 0.855 0.76 0.855 0.54 0.935 0.54 ;
  END
END SPDFF2RX2

MACRO SPDFF4RX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SPDFF4RX1 0 0 ;
  SIZE 20.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.83755 LAYER Metal1 ;
    ANTENNADIFFAREA 21.9111 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8982 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.17919175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 97.83567125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.84 1.11 5.71 1.11 5.71 0.96 5.66 0.96 5.66 0.76 5.725 0.76 5.725 0.6 5.73 0.6 5.73 0.54 5.805 0.54 5.805 1.05 5.84 1.05 ;
    END
  END Q2
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.83755 LAYER Metal1 ;
    ANTENNADIFFAREA 16.969525 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8982 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.17919175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 97.83567125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.19 1.11 5.06 1.11 5.06 0.54 5.155 0.54 5.155 1.05 5.19 1.05 ;
    END
  END Q2N
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.785 0.775 8.74 0.775 8.74 0.875 8.66 0.875 8.66 0.62 8.785 0.62 ;
    END
  END D2
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.429625 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1296 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.031057 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 104.56018525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.735 1.35 17.735 1.35 17.735 1.375 17.335 1.375 17.335 1.35 12.735 1.35 12.735 1.375 12.335 1.375 12.335 1.35 10.755 1.35 10.755 1.465 10.46 1.465 10.46 1.35 8.465 1.35 8.465 1.375 8.065 1.375 8.065 1.35 3.465 1.35 3.465 1.375 3.065 1.375 3.065 1.35 0.065 1.35 0.065 1.29 3.125 1.29 3.125 1.315 3.41 1.315 3.41 1.29 8.125 1.29 8.125 1.315 8.41 1.315 8.41 1.29 12.39 1.29 12.39 1.315 12.675 1.315 12.675 1.29 17.39 1.29 17.39 1.315 17.675 1.315 17.675 1.29 20.735 1.29 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1296 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 59.1435185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.735 0.41 16.57 0.41 16.57 0.7 16.835 0.7 16.835 0.865 16.775 0.865 16.775 0.76 16.51 0.76 16.51 0.41 16.145 0.41 16.145 0.895 16.06 0.895 16.06 0.41 11.57 0.41 11.57 0.7 11.835 0.7 11.835 0.865 11.775 0.865 11.775 0.76 11.51 0.76 11.51 0.41 11.145 0.41 11.145 0.895 11.06 0.895 11.06 0.41 9.74 0.41 9.74 0.895 9.655 0.895 9.655 0.41 9.29 0.41 9.29 0.76 9.025 0.76 9.025 0.865 8.965 0.865 8.965 0.7 9.23 0.7 9.23 0.41 4.74 0.41 4.74 0.895 4.655 0.895 4.655 0.41 4.29 0.41 4.29 0.76 4.025 0.76 4.025 0.865 3.965 0.865 3.965 0.7 4.23 0.7 4.23 0.41 0.065 0.41 0.065 0.35 20.735 0.35 ;
    END
  END SE
  PIN SI2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 9.39 0.625 9.565 0.77 ;
    END
  END SI2
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.83755 LAYER Metal1 ;
    ANTENNADIFFAREA 18.759525 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8982 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.17919175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 97.83567125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.84 1.11 0.71 1.11 0.71 0.96 0.66 0.96 0.66 0.76 0.725 0.76 0.725 0.6 0.73 0.6 0.73 0.54 0.805 0.54 0.805 1.05 0.84 1.05 ;
    END
  END Q1
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.83755 LAYER Metal1 ;
    ANTENNADIFFAREA 16.969525 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8982 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.17919175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 97.83567125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.19 1.11 0.06 1.11 0.06 0.54 0.155 0.54 0.155 1.05 0.19 1.05 ;
    END
  END Q1N
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.785 0.775 3.74 0.775 3.74 0.875 3.66 0.875 3.66 0.62 3.785 0.62 ;
    END
  END D1
  PIN SI1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.39 0.625 4.565 0.77 ;
    END
  END SI1
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.445 0.77 10.625 0.92 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.8 1.77 0 1.77 0 1.65 0.3 1.65 0.3 1.54 0.42 1.54 0.42 1.65 0.955 1.65 0.955 1.54 1.075 1.54 1.075 1.65 1.53 1.65 1.53 1.54 1.65 1.54 1.65 1.65 2.445 1.65 2.445 1.54 2.565 1.54 2.565 1.65 2.795 1.65 2.795 1.54 2.915 1.54 2.915 1.65 3.675 1.65 3.675 1.54 3.795 1.54 3.795 1.65 4.465 1.65 4.465 1.54 4.585 1.54 4.585 1.65 5.3 1.65 5.3 1.54 5.42 1.54 5.42 1.65 5.955 1.65 5.955 1.54 6.075 1.54 6.075 1.65 6.53 1.65 6.53 1.54 6.65 1.54 6.65 1.65 7.445 1.65 7.445 1.54 7.565 1.54 7.565 1.65 7.795 1.65 7.795 1.54 7.915 1.54 7.915 1.65 8.675 1.65 8.675 1.54 8.795 1.54 8.795 1.65 9.465 1.65 9.465 1.54 9.585 1.54 9.585 1.65 10.33 1.65 10.33 1.54 10.45 1.54 10.45 1.65 11.215 1.65 11.215 1.54 11.335 1.54 11.335 1.65 12.005 1.65 12.005 1.54 12.125 1.54 12.125 1.65 12.885 1.65 12.885 1.54 13.005 1.54 13.005 1.65 13.235 1.65 13.235 1.54 13.355 1.54 13.355 1.65 14.15 1.65 14.15 1.54 14.27 1.54 14.27 1.65 14.725 1.65 14.725 1.54 14.845 1.54 14.845 1.65 15.38 1.65 15.38 1.54 15.5 1.54 15.5 1.65 16.215 1.65 16.215 1.54 16.335 1.54 16.335 1.65 17.005 1.65 17.005 1.54 17.125 1.54 17.125 1.65 17.885 1.65 17.885 1.54 18.005 1.54 18.005 1.65 18.235 1.65 18.235 1.54 18.355 1.54 18.355 1.65 19.15 1.65 19.15 1.54 19.27 1.54 19.27 1.65 19.725 1.65 19.725 1.54 19.845 1.54 19.845 1.65 20.38 1.65 20.38 1.54 20.5 1.54 20.5 1.65 20.8 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.8 0.06 20.5 0.06 20.5 0.17 20.38 0.17 20.38 0.06 19.895 0.06 19.895 0.17 19.775 0.17 19.775 0.06 19.27 0.06 19.27 0.17 19.15 0.17 19.15 0.06 18.255 0.06 18.255 0.17 18.135 0.17 18.135 0.06 17.15 0.06 17.15 0.17 17.03 0.17 17.03 0.06 16.335 0.06 16.335 0.17 16.215 0.17 16.215 0.06 15.5 0.06 15.5 0.17 15.38 0.17 15.38 0.06 14.895 0.06 14.895 0.17 14.775 0.17 14.775 0.06 14.27 0.06 14.27 0.17 14.15 0.17 14.15 0.06 13.255 0.06 13.255 0.17 13.135 0.17 13.135 0.06 12.15 0.06 12.15 0.17 12.03 0.17 12.03 0.06 11.335 0.06 11.335 0.17 11.215 0.17 11.215 0.06 10.45 0.06 10.45 0.17 10.325 0.17 10.325 0.06 9.585 0.06 9.585 0.17 9.465 0.17 9.465 0.06 8.77 0.06 8.77 0.17 8.65 0.17 8.65 0.06 7.665 0.06 7.665 0.17 7.545 0.17 7.545 0.06 6.65 0.06 6.65 0.17 6.53 0.17 6.53 0.06 6.025 0.06 6.025 0.17 5.905 0.17 5.905 0.06 5.42 0.06 5.42 0.17 5.3 0.17 5.3 0.06 4.585 0.06 4.585 0.17 4.465 0.17 4.465 0.06 3.77 0.06 3.77 0.17 3.65 0.17 3.65 0.06 2.665 0.06 2.665 0.17 2.545 0.17 2.545 0.06 1.65 0.06 1.65 0.17 1.53 0.17 1.53 0.06 1.025 0.06 1.025 0.17 0.905 0.17 0.905 0.06 0.42 0.06 0.42 0.17 0.3 0.17 0.3 0.06 0 0.06 0 -0.06 20.8 -0.06 ;
    END
  END VSS
  PIN Q4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.83755 LAYER Metal1 ;
    ANTENNADIFFAREA 25.88645 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8982 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.17919175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 97.83567125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.14 0.96 20.09 0.96 20.09 1.11 19.96 1.11 19.96 1.05 19.995 1.05 19.995 0.54 20.07 0.54 20.07 0.6 20.075 0.6 20.075 0.76 20.14 0.76 ;
    END
  END Q4
  PIN Q4N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.83755 LAYER Metal1 ;
    ANTENNADIFFAREA 25.205025 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8982 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.17919175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 97.83567125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 20.74 1.11 20.61 1.11 20.61 1.05 20.645 1.05 20.645 0.54 20.74 0.54 ;
    END
  END Q4N
  PIN D4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 17.14 0.875 17.06 0.875 17.06 0.775 17.015 0.775 17.015 0.62 17.14 0.62 ;
    END
  END D4
  PIN SI4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 16.235 0.625 16.41 0.77 ;
    END
  END SI4
  PIN Q3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.83755 LAYER Metal1 ;
    ANTENNADIFFAREA 22.024725 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8982 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.17919175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 97.83567125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.14 0.96 15.09 0.96 15.09 1.11 14.96 1.11 14.96 1.05 14.995 1.05 14.995 0.54 15.07 0.54 15.07 0.6 15.075 0.6 15.075 0.76 15.14 0.76 ;
    END
  END Q3
  PIN Q3N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.83755 LAYER Metal1 ;
    ANTENNADIFFAREA 23.929175 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.8982 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.17919175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 97.83567125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 15.74 1.11 15.61 1.11 15.61 1.05 15.645 1.05 15.645 0.54 15.74 0.54 ;
    END
  END Q3N
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 12.14 0.875 12.06 0.875 12.06 0.775 12.015 0.775 12.015 0.62 12.14 0.62 ;
    END
  END D3
  PIN SI3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.235 0.625 11.41 0.77 ;
    END
  END SI3
  OBS
    LAYER Metal1 ;
      POLYGON 20.735 0.29 0.065 0.29 0.065 0.23 4.66 0.23 4.66 0.205 4.8 0.205 4.8 0.23 9.66 0.23 9.66 0.205 9.8 0.205 9.8 0.23 11 0.23 11 0.205 11.14 0.205 11.14 0.23 16 0.23 16 0.205 16.14 0.205 16.14 0.23 20.735 0.23 ;
      POLYGON 20.735 1.23 17.615 1.23 17.615 1.255 17.45 1.255 17.45 1.23 12.615 1.23 12.615 1.255 12.45 1.255 12.45 1.23 8.35 1.23 8.35 1.255 8.185 1.255 8.185 1.23 3.35 1.23 3.35 1.255 3.185 1.255 3.185 1.23 0.065 1.23 0.065 1.17 1.835 1.17 1.835 0.665 1.895 0.665 1.895 1.17 2.165 1.17 2.165 0.865 2.105 0.865 2.105 0.805 2.225 0.805 2.225 1.17 4.64 1.17 4.64 1.15 4.78 1.15 4.78 1.17 6.835 1.17 6.835 0.665 6.895 0.665 6.895 1.17 7.165 1.17 7.165 0.865 7.105 0.865 7.105 0.805 7.225 0.805 7.225 1.17 9.64 1.17 9.64 1.15 9.78 1.15 9.78 1.17 10.3 1.17 10.3 0.895 10.26 0.895 10.26 0.495 10.36 0.495 10.36 0.625 10.565 0.625 10.565 0.505 10.625 0.505 10.625 0.705 10.36 0.705 10.36 1.005 10.655 1.005 10.655 1.065 10.36 1.065 10.36 1.17 11.02 1.17 11.02 1.15 11.16 1.15 11.16 1.17 13.575 1.17 13.575 0.805 13.695 0.805 13.695 0.865 13.635 0.865 13.635 1.17 13.905 1.17 13.905 0.665 13.965 0.665 13.965 1.17 16.02 1.17 16.02 1.15 16.16 1.15 16.16 1.17 18.575 1.17 18.575 0.805 18.695 0.805 18.695 0.865 18.635 0.865 18.635 1.17 18.905 1.17 18.905 0.665 18.965 0.665 18.965 1.17 20.735 1.17 ;
      POLYGON 20.73 1.48 17.84 1.48 17.84 1.495 17.22 1.495 17.22 1.48 17.005 1.48 17.005 1.42 17.275 1.42 17.275 1.435 17.78 1.435 17.78 1.42 20.73 1.42 ;
      POLYGON 20.545 0.84 20.29 0.84 20.29 1.02 20.21 1.02 20.21 0.54 20.29 0.54 20.29 0.76 20.545 0.76 ;
      POLYGON 19.925 0.82 19.645 0.82 19.645 1.1 19.075 1.1 19.075 0.68 19.135 0.68 19.135 1.04 19.585 1.04 19.585 0.485 19.645 0.485 19.645 0.76 19.925 0.76 ;
      POLYGON 19.515 0.825 19.455 0.825 19.455 0.66 19.4 0.66 19.4 0.575 18.82 0.575 18.82 1.055 18.76 1.055 18.76 0.575 18.71 0.575 18.71 0.495 19.46 0.495 19.46 0.6 19.515 0.6 ;
      RECT 19.235 0.735 19.395 0.96 ;
      POLYGON 18.54 0.575 18.51 0.575 18.51 1.055 18.45 1.055 18.45 0.74 17.855 0.74 17.855 0.68 18.45 0.68 18.45 0.575 18.42 0.575 18.42 0.515 18.54 0.515 ;
      POLYGON 18.37 0.86 17.52 0.86 17.52 1.045 17.46 1.045 17.46 0.8 17.645 0.8 17.645 0.575 17.61 0.575 17.61 0.515 17.74 0.515 17.74 0.575 17.705 0.575 17.705 0.8 18.37 0.8 ;
      RECT 17.635 0.95 18.135 1.03 ;
      POLYGON 17.53 0.575 17.5 0.575 17.5 0.73 17.4 0.73 17.4 0.95 17.315 0.95 17.315 1.065 16.615 1.065 16.615 1.005 16.895 1.005 16.895 0.54 16.655 0.54 16.655 0.48 16.955 0.48 16.955 1.005 17.255 1.005 17.255 0.89 17.34 0.89 17.34 0.67 17.44 0.67 17.44 0.575 17.41 0.575 17.41 0.515 17.53 0.515 ;
      POLYGON 16.67 0.905 16.315 0.905 16.315 1.065 15.925 1.065 15.925 0.51 15.985 0.51 15.985 1.005 16.255 1.005 16.255 0.845 16.67 0.845 ;
      POLYGON 16.495 1.48 12.84 1.48 12.84 1.495 12.22 1.495 12.22 1.48 12.005 1.48 12.005 1.42 12.275 1.42 12.275 1.435 12.78 1.435 12.78 1.42 16.495 1.42 ;
      POLYGON 15.545 0.84 15.29 0.84 15.29 1.02 15.21 1.02 15.21 0.54 15.29 0.54 15.29 0.76 15.545 0.76 ;
      POLYGON 14.925 0.82 14.645 0.82 14.645 1.1 14.075 1.1 14.075 0.68 14.135 0.68 14.135 1.04 14.585 1.04 14.585 0.485 14.645 0.485 14.645 0.76 14.925 0.76 ;
      POLYGON 14.515 0.825 14.455 0.825 14.455 0.66 14.4 0.66 14.4 0.575 13.82 0.575 13.82 1.055 13.76 1.055 13.76 0.575 13.71 0.575 13.71 0.495 14.46 0.495 14.46 0.6 14.515 0.6 ;
      RECT 14.235 0.735 14.395 0.96 ;
      POLYGON 13.54 0.575 13.51 0.575 13.51 1.055 13.45 1.055 13.45 0.74 12.855 0.74 12.855 0.68 13.45 0.68 13.45 0.575 13.42 0.575 13.42 0.515 13.54 0.515 ;
      POLYGON 13.37 0.86 12.52 0.86 12.52 1.045 12.46 1.045 12.46 0.8 12.645 0.8 12.645 0.575 12.61 0.575 12.61 0.515 12.74 0.515 12.74 0.575 12.705 0.575 12.705 0.8 13.37 0.8 ;
      RECT 12.635 0.95 13.135 1.03 ;
      POLYGON 12.53 0.575 12.5 0.575 12.5 0.73 12.4 0.73 12.4 0.95 12.315 0.95 12.315 1.065 11.615 1.065 11.615 1.005 11.895 1.005 11.895 0.54 11.655 0.54 11.655 0.48 11.955 0.48 11.955 1.005 12.255 1.005 12.255 0.89 12.34 0.89 12.34 0.67 12.44 0.67 12.44 0.575 12.41 0.575 12.41 0.515 12.53 0.515 ;
      POLYGON 11.67 0.905 11.315 0.905 11.315 1.065 10.925 1.065 10.925 0.51 10.985 0.51 10.985 1.005 11.255 1.005 11.255 0.845 11.67 0.845 ;
      RECT 10.925 1.42 11.495 1.48 ;
      POLYGON 10.2 1.1 10.06 1.1 10.06 0.77 10.14 0.77 10.14 0.495 10.2 0.495 ;
      POLYGON 9.875 1.065 9.485 1.065 9.485 0.905 9.13 0.905 9.13 0.845 9.545 0.845 9.545 1.005 9.815 1.005 9.815 0.51 9.875 0.51 ;
      RECT 9.305 1.42 9.875 1.48 ;
      POLYGON 9.185 1.065 8.485 1.065 8.485 0.95 8.4 0.95 8.4 0.73 8.3 0.73 8.3 0.575 8.27 0.575 8.27 0.515 8.39 0.515 8.39 0.575 8.36 0.575 8.36 0.67 8.46 0.67 8.46 0.89 8.545 0.89 8.545 1.005 8.845 1.005 8.845 0.48 9.145 0.48 9.145 0.54 8.905 0.54 8.905 1.005 9.185 1.005 ;
      POLYGON 8.795 1.48 8.58 1.48 8.58 1.495 7.96 1.495 7.96 1.48 4.305 1.48 4.305 1.42 8.02 1.42 8.02 1.435 8.525 1.435 8.525 1.42 8.795 1.42 ;
      POLYGON 8.34 1.045 8.28 1.045 8.28 0.86 7.43 0.86 7.43 0.8 8.095 0.8 8.095 0.575 8.06 0.575 8.06 0.515 8.19 0.515 8.19 0.575 8.155 0.575 8.155 0.8 8.34 0.8 ;
      RECT 7.665 0.95 8.165 1.03 ;
      POLYGON 7.945 0.74 7.35 0.74 7.35 1.055 7.29 1.055 7.29 0.575 7.26 0.575 7.26 0.515 7.38 0.515 7.38 0.575 7.35 0.575 7.35 0.68 7.945 0.68 ;
      POLYGON 7.09 0.575 7.04 0.575 7.04 1.055 6.98 1.055 6.98 0.575 6.4 0.575 6.4 0.66 6.345 0.66 6.345 0.825 6.285 0.825 6.285 0.6 6.34 0.6 6.34 0.495 7.09 0.495 ;
      POLYGON 6.725 1.1 6.155 1.1 6.155 0.82 5.875 0.82 5.875 0.76 6.155 0.76 6.155 0.485 6.215 0.485 6.215 1.04 6.665 1.04 6.665 0.68 6.725 0.68 ;
      RECT 6.405 0.735 6.565 0.96 ;
      POLYGON 5.59 1.02 5.51 1.02 5.51 0.84 5.255 0.84 5.255 0.76 5.51 0.76 5.51 0.54 5.59 0.54 ;
      POLYGON 4.875 1.065 4.485 1.065 4.485 0.905 4.13 0.905 4.13 0.845 4.545 0.845 4.545 1.005 4.815 1.005 4.815 0.51 4.875 0.51 ;
      POLYGON 4.185 1.065 3.485 1.065 3.485 0.95 3.4 0.95 3.4 0.73 3.3 0.73 3.3 0.575 3.27 0.575 3.27 0.515 3.39 0.515 3.39 0.575 3.36 0.575 3.36 0.67 3.46 0.67 3.46 0.89 3.545 0.89 3.545 1.005 3.845 1.005 3.845 0.48 4.145 0.48 4.145 0.54 3.905 0.54 3.905 1.005 4.185 1.005 ;
      POLYGON 3.795 1.48 3.58 1.48 3.58 1.495 2.96 1.495 2.96 1.48 0.07 1.48 0.07 1.42 3.02 1.42 3.02 1.435 3.525 1.435 3.525 1.42 3.795 1.42 ;
      POLYGON 3.34 1.045 3.28 1.045 3.28 0.86 2.43 0.86 2.43 0.8 3.095 0.8 3.095 0.575 3.06 0.575 3.06 0.515 3.19 0.515 3.19 0.575 3.155 0.575 3.155 0.8 3.34 0.8 ;
      RECT 2.665 0.95 3.165 1.03 ;
      POLYGON 2.945 0.74 2.35 0.74 2.35 1.055 2.29 1.055 2.29 0.575 2.26 0.575 2.26 0.515 2.38 0.515 2.38 0.575 2.35 0.575 2.35 0.68 2.945 0.68 ;
      POLYGON 2.09 0.575 2.04 0.575 2.04 1.055 1.98 1.055 1.98 0.575 1.4 0.575 1.4 0.66 1.345 0.66 1.345 0.825 1.285 0.825 1.285 0.6 1.34 0.6 1.34 0.495 2.09 0.495 ;
      POLYGON 1.725 1.1 1.155 1.1 1.155 0.82 0.875 0.82 0.875 0.76 1.155 0.76 1.155 0.485 1.215 0.485 1.215 1.04 1.665 1.04 1.665 0.68 1.725 0.68 ;
      RECT 1.405 0.735 1.565 0.96 ;
      POLYGON 0.59 1.02 0.51 1.02 0.51 0.84 0.255 0.84 0.255 0.76 0.51 0.76 0.51 0.54 0.59 0.54 ;
  END
END SPDFF4RX1

MACRO SPDFF4RX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SPDFF4RX2 0 0 ;
  SIZE 23.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.71595 LAYER Metal1 ;
    ANTENNADIFFAREA 19.511475 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.1601 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.961081 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 78.241531 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.86 0.54 7.015 1.11 ;
    END
  END Q2
  PIN D2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.985 0.775 9.94 0.775 9.94 0.875 9.86 0.875 9.86 0.62 9.985 0.62 ;
    END
  END D2
  PIN Q2N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.71595 LAYER Metal1 ;
    ANTENNADIFFAREA 19.14045 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.1601 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.961081 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 78.241531 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.005 0.54 6.145 1.11 ;
    END
  END Q2N
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.373875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1575 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.72301575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 82.5714285 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 21.48 1.35 19.535 1.35 19.535 1.375 19.135 1.375 19.135 1.35 13.935 1.35 13.935 1.375 13.535 1.375 13.535 1.35 11.945 1.35 11.945 1.465 11.66 1.465 11.66 1.35 9.665 1.35 9.665 1.375 9.265 1.375 9.265 1.35 4.065 1.35 4.065 1.375 3.665 1.375 3.665 1.35 1.72 1.35 1.72 1.29 3.725 1.29 3.725 1.315 4.01 1.315 4.01 1.29 9.325 1.29 9.325 1.315 9.61 1.315 9.61 1.29 13.59 1.29 13.59 1.315 13.875 1.315 13.875 1.29 19.19 1.29 19.19 1.315 19.475 1.315 19.475 1.29 21.48 1.29 ;
    END
  END RN
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1296 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 57.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 21.48 0.41 18.37 0.41 18.37 0.7 18.635 0.7 18.635 0.865 18.575 0.865 18.575 0.76 18.31 0.76 18.31 0.41 17.945 0.41 17.945 0.895 17.86 0.895 17.86 0.41 12.77 0.41 12.77 0.7 13.035 0.7 13.035 0.865 12.975 0.865 12.975 0.76 12.71 0.76 12.71 0.41 12.345 0.41 12.345 0.895 12.26 0.895 12.26 0.41 10.94 0.41 10.94 0.895 10.855 0.895 10.855 0.41 10.49 0.41 10.49 0.76 10.225 0.76 10.225 0.865 10.165 0.865 10.165 0.7 10.43 0.7 10.43 0.41 5.34 0.41 5.34 0.895 5.255 0.895 5.255 0.41 4.89 0.41 4.89 0.76 4.625 0.76 4.625 0.865 4.565 0.865 4.565 0.7 4.83 0.7 4.83 0.41 1.72 0.41 1.72 0.35 21.48 0.35 ;
    END
  END SE
  PIN SI2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 10.59 0.625 10.765 0.77 ;
    END
  END SI2
  PIN Q1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.71595 LAYER Metal1 ;
    ANTENNADIFFAREA 22.377125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.1601 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.961081 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 78.241531 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.26 0.54 1.415 1.11 ;
    END
  END Q1
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.385 0.775 4.34 0.775 4.34 0.875 4.26 0.875 4.26 0.62 4.385 0.62 ;
    END
  END D1
  PIN Q1N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.71595 LAYER Metal1 ;
    ANTENNADIFFAREA 20.422525 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.1601 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.961081 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 78.241531 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.405 0.54 0.545 1.11 ;
    END
  END Q1N
  PIN SI1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.99 0.625 5.165 0.77 ;
    END
  END SI1
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 11.645 0.77 11.825 0.92 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.2 1.77 0 1.77 0 1.65 0.24 1.65 0.24 1.54 0.36 1.54 0.36 1.65 0.61 1.65 0.61 1.54 0.765 1.54 0.765 1.65 1.065 1.65 1.065 1.54 1.185 1.54 1.185 1.65 1.555 1.65 1.555 1.54 1.675 1.54 1.675 1.65 2.13 1.65 2.13 1.54 2.25 1.54 2.25 1.65 3.045 1.65 3.045 1.54 3.165 1.54 3.165 1.65 3.395 1.65 3.395 1.54 3.515 1.54 3.515 1.65 4.275 1.65 4.275 1.54 4.395 1.54 4.395 1.65 5.065 1.65 5.065 1.54 5.185 1.54 5.185 1.65 5.84 1.65 5.84 1.54 5.96 1.54 5.96 1.65 6.21 1.65 6.21 1.54 6.365 1.54 6.365 1.65 6.665 1.65 6.665 1.54 6.785 1.54 6.785 1.65 7.155 1.65 7.155 1.54 7.275 1.54 7.275 1.65 7.73 1.65 7.73 1.54 7.85 1.54 7.85 1.65 8.645 1.65 8.645 1.54 8.765 1.54 8.765 1.65 8.995 1.65 8.995 1.54 9.115 1.54 9.115 1.65 9.875 1.65 9.875 1.54 9.995 1.54 9.995 1.65 10.665 1.65 10.665 1.54 10.785 1.54 10.785 1.65 11.53 1.65 11.53 1.54 11.65 1.54 11.65 1.65 12.415 1.65 12.415 1.54 12.535 1.54 12.535 1.65 13.205 1.65 13.205 1.54 13.325 1.54 13.325 1.65 14.085 1.65 14.085 1.54 14.205 1.54 14.205 1.65 14.435 1.65 14.435 1.54 14.555 1.54 14.555 1.65 15.35 1.65 15.35 1.54 15.47 1.54 15.47 1.65 15.925 1.65 15.925 1.54 16.045 1.54 16.045 1.65 16.415 1.65 16.415 1.54 16.535 1.54 16.535 1.65 16.835 1.65 16.835 1.54 16.99 1.54 16.99 1.65 17.24 1.65 17.24 1.54 17.36 1.54 17.36 1.65 18.015 1.65 18.015 1.54 18.135 1.54 18.135 1.65 18.805 1.65 18.805 1.54 18.925 1.54 18.925 1.65 19.685 1.65 19.685 1.54 19.805 1.54 19.805 1.65 20.035 1.65 20.035 1.54 20.155 1.54 20.155 1.65 20.95 1.65 20.95 1.54 21.07 1.54 21.07 1.65 21.525 1.65 21.525 1.54 21.645 1.54 21.645 1.65 22.015 1.65 22.015 1.54 22.135 1.54 22.135 1.65 22.435 1.65 22.435 1.54 22.59 1.54 22.59 1.65 22.84 1.65 22.84 1.54 22.96 1.54 22.96 1.65 23.2 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 23.2 0.06 22.96 0.06 22.96 0.17 22.84 0.17 22.84 0.06 22.59 0.06 22.59 0.17 22.47 0.17 22.47 0.06 22.135 0.06 22.135 0.17 22.015 0.17 22.015 0.06 21.695 0.06 21.695 0.17 21.575 0.17 21.575 0.06 21.07 0.06 21.07 0.17 20.95 0.17 20.95 0.06 20.055 0.06 20.055 0.17 19.935 0.17 19.935 0.06 18.95 0.06 18.95 0.17 18.83 0.17 18.83 0.06 18.135 0.06 18.135 0.17 18.015 0.17 18.015 0.06 17.36 0.06 17.36 0.17 17.24 0.17 17.24 0.06 16.99 0.06 16.99 0.17 16.87 0.17 16.87 0.06 16.535 0.06 16.535 0.17 16.415 0.17 16.415 0.06 16.095 0.06 16.095 0.17 15.975 0.17 15.975 0.06 15.47 0.06 15.47 0.17 15.35 0.17 15.35 0.06 14.455 0.06 14.455 0.17 14.335 0.17 14.335 0.06 13.35 0.06 13.35 0.17 13.23 0.17 13.23 0.06 12.535 0.06 12.535 0.17 12.415 0.17 12.415 0.06 11.65 0.06 11.65 0.17 11.525 0.17 11.525 0.06 10.785 0.06 10.785 0.17 10.665 0.17 10.665 0.06 9.97 0.06 9.97 0.17 9.85 0.17 9.85 0.06 8.865 0.06 8.865 0.17 8.745 0.17 8.745 0.06 7.85 0.06 7.85 0.17 7.73 0.17 7.73 0.06 7.225 0.06 7.225 0.17 7.105 0.17 7.105 0.06 6.785 0.06 6.785 0.17 6.665 0.17 6.665 0.06 6.33 0.06 6.33 0.17 6.21 0.17 6.21 0.06 5.96 0.06 5.96 0.17 5.84 0.17 5.84 0.06 5.185 0.06 5.185 0.17 5.065 0.17 5.065 0.06 4.37 0.06 4.37 0.17 4.25 0.17 4.25 0.06 3.265 0.06 3.265 0.17 3.145 0.17 3.145 0.06 2.25 0.06 2.25 0.17 2.13 0.17 2.13 0.06 1.625 0.06 1.625 0.17 1.505 0.17 1.505 0.06 1.185 0.06 1.185 0.17 1.065 0.17 1.065 0.06 0.73 0.06 0.73 0.17 0.61 0.17 0.61 0.06 0.36 0.06 0.36 0.17 0.24 0.17 0.24 0.06 0 0.06 0 -0.06 23.2 -0.06 ;
    END
  END VSS
  PIN Q4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.71595 LAYER Metal1 ;
    ANTENNADIFFAREA 30.152275 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.1601 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.961081 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 78.241531 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 21.785 0.54 21.94 1.11 ;
    END
  END Q4
  PIN D4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 18.94 0.875 18.86 0.875 18.86 0.775 18.815 0.775 18.815 0.62 18.94 0.62 ;
    END
  END D4
  PIN Q4N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.71595 LAYER Metal1 ;
    ANTENNADIFFAREA 29.839075 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.1601 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.961081 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 78.241531 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 22.655 0.54 22.795 1.11 ;
    END
  END Q4N
  PIN SI4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 18.035 0.625 18.21 0.77 ;
    END
  END SI4
  PIN Q3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.71595 LAYER Metal1 ;
    ANTENNADIFFAREA 24.068275 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.1601 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.961081 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 78.241531 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 16.185 0.54 16.34 1.11 ;
    END
  END Q3
  PIN D3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 13.34 0.875 13.26 0.875 13.26 0.775 13.215 0.775 13.215 0.62 13.34 0.62 ;
    END
  END D3
  PIN Q3N
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.71595 LAYER Metal1 ;
    ANTENNADIFFAREA 23.755075 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.1601 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.961081 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 78.241531 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 17.055 0.54 17.195 1.11 ;
    END
  END Q3N
  PIN SI3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 12.435 0.625 12.61 0.77 ;
    END
  END SI3
  OBS
    LAYER Metal1 ;
      POLYGON 22.57 0.85 22.51 0.85 22.51 0.82 22.345 0.82 22.345 1.02 22.265 1.02 22.265 0.54 22.345 0.54 22.345 0.76 22.51 0.76 22.51 0.725 22.57 0.725 ;
      POLYGON 21.725 0.82 21.445 0.82 21.445 1.1 20.875 1.1 20.875 0.68 20.935 0.68 20.935 1.04 21.385 1.04 21.385 0.485 21.445 0.485 21.445 0.76 21.725 0.76 ;
      POLYGON 21.48 0.29 1.72 0.29 1.72 0.23 5.26 0.23 5.26 0.205 5.4 0.205 5.4 0.23 10.86 0.23 10.86 0.205 11 0.205 11 0.23 12.2 0.23 12.2 0.205 12.34 0.205 12.34 0.23 17.8 0.23 17.8 0.205 17.94 0.205 17.94 0.23 21.48 0.23 ;
      POLYGON 21.48 1.23 19.415 1.23 19.415 1.255 19.25 1.255 19.25 1.23 13.815 1.23 13.815 1.255 13.65 1.255 13.65 1.23 9.55 1.23 9.55 1.255 9.385 1.255 9.385 1.23 3.95 1.23 3.95 1.255 3.785 1.255 3.785 1.23 1.72 1.23 1.72 1.17 2.435 1.17 2.435 0.665 2.495 0.665 2.495 1.17 2.765 1.17 2.765 0.865 2.705 0.865 2.705 0.805 2.825 0.805 2.825 1.17 5.24 1.17 5.24 1.15 5.38 1.15 5.38 1.17 8.035 1.17 8.035 0.665 8.095 0.665 8.095 1.17 8.365 1.17 8.365 0.865 8.305 0.865 8.305 0.805 8.425 0.805 8.425 1.17 10.84 1.17 10.84 1.15 10.98 1.15 10.98 1.17 11.5 1.17 11.5 0.895 11.46 0.895 11.46 0.495 11.56 0.495 11.56 0.625 11.765 0.625 11.765 0.505 11.825 0.505 11.825 0.705 11.56 0.705 11.56 1.005 11.855 1.005 11.855 1.065 11.56 1.065 11.56 1.17 12.22 1.17 12.22 1.15 12.36 1.15 12.36 1.17 14.775 1.17 14.775 0.805 14.895 0.805 14.895 0.865 14.835 0.865 14.835 1.17 15.105 1.17 15.105 0.665 15.165 0.665 15.165 1.17 17.82 1.17 17.82 1.15 17.96 1.15 17.96 1.17 20.375 1.17 20.375 0.805 20.495 0.805 20.495 0.865 20.435 0.865 20.435 1.17 20.705 1.17 20.705 0.665 20.765 0.665 20.765 1.17 21.48 1.17 ;
      POLYGON 21.475 1.48 19.64 1.48 19.64 1.495 19.02 1.495 19.02 1.48 18.805 1.48 18.805 1.42 19.075 1.42 19.075 1.435 19.58 1.435 19.58 1.42 21.475 1.42 ;
      POLYGON 21.315 0.825 21.255 0.825 21.255 0.66 21.2 0.66 21.2 0.575 20.62 0.575 20.62 1.055 20.56 1.055 20.56 0.575 20.51 0.575 20.51 0.495 21.26 0.495 21.26 0.6 21.315 0.6 ;
      RECT 21.035 0.735 21.195 0.96 ;
      POLYGON 20.34 0.575 20.31 0.575 20.31 1.055 20.25 1.055 20.25 0.74 19.655 0.74 19.655 0.68 20.25 0.68 20.25 0.575 20.22 0.575 20.22 0.515 20.34 0.515 ;
      POLYGON 20.17 0.86 19.32 0.86 19.32 1.045 19.26 1.045 19.26 0.8 19.445 0.8 19.445 0.575 19.41 0.575 19.41 0.515 19.54 0.515 19.54 0.575 19.505 0.575 19.505 0.8 20.17 0.8 ;
      RECT 19.435 0.95 19.935 1.03 ;
      POLYGON 19.33 0.575 19.3 0.575 19.3 0.73 19.2 0.73 19.2 0.95 19.115 0.95 19.115 1.065 18.415 1.065 18.415 1.005 18.695 1.005 18.695 0.54 18.455 0.54 18.455 0.48 18.755 0.48 18.755 1.005 19.055 1.005 19.055 0.89 19.14 0.89 19.14 0.67 19.24 0.67 19.24 0.575 19.21 0.575 19.21 0.515 19.33 0.515 ;
      POLYGON 18.47 0.905 18.115 0.905 18.115 1.065 17.725 1.065 17.725 0.51 17.785 0.51 17.785 1.005 18.055 1.005 18.055 0.845 18.47 0.845 ;
      POLYGON 18.295 1.48 14.04 1.48 14.04 1.495 13.42 1.495 13.42 1.48 13.205 1.48 13.205 1.42 13.475 1.42 13.475 1.435 13.98 1.435 13.98 1.42 18.295 1.42 ;
      POLYGON 16.97 0.85 16.91 0.85 16.91 0.82 16.745 0.82 16.745 1.02 16.665 1.02 16.665 0.54 16.745 0.54 16.745 0.76 16.91 0.76 16.91 0.725 16.97 0.725 ;
      POLYGON 16.125 0.82 15.845 0.82 15.845 1.1 15.275 1.1 15.275 0.68 15.335 0.68 15.335 1.04 15.785 1.04 15.785 0.485 15.845 0.485 15.845 0.76 16.125 0.76 ;
      POLYGON 15.715 0.825 15.655 0.825 15.655 0.66 15.6 0.66 15.6 0.575 15.02 0.575 15.02 1.055 14.96 1.055 14.96 0.575 14.91 0.575 14.91 0.495 15.66 0.495 15.66 0.6 15.715 0.6 ;
      RECT 15.435 0.735 15.595 0.96 ;
      POLYGON 14.74 0.575 14.71 0.575 14.71 1.055 14.65 1.055 14.65 0.74 14.055 0.74 14.055 0.68 14.65 0.68 14.65 0.575 14.62 0.575 14.62 0.515 14.74 0.515 ;
      POLYGON 14.57 0.86 13.72 0.86 13.72 1.045 13.66 1.045 13.66 0.8 13.845 0.8 13.845 0.575 13.81 0.575 13.81 0.515 13.94 0.515 13.94 0.575 13.905 0.575 13.905 0.8 14.57 0.8 ;
      RECT 13.835 0.95 14.335 1.03 ;
      POLYGON 13.73 0.575 13.7 0.575 13.7 0.73 13.6 0.73 13.6 0.95 13.515 0.95 13.515 1.065 12.815 1.065 12.815 1.005 13.095 1.005 13.095 0.54 12.855 0.54 12.855 0.48 13.155 0.48 13.155 1.005 13.455 1.005 13.455 0.89 13.54 0.89 13.54 0.67 13.64 0.67 13.64 0.575 13.61 0.575 13.61 0.515 13.73 0.515 ;
      POLYGON 12.87 0.905 12.515 0.905 12.515 1.065 12.125 1.065 12.125 0.51 12.185 0.51 12.185 1.005 12.455 1.005 12.455 0.845 12.87 0.845 ;
      RECT 12.125 1.42 12.695 1.48 ;
      POLYGON 11.4 1.1 11.26 1.1 11.26 0.77 11.34 0.77 11.34 0.495 11.4 0.495 ;
      POLYGON 11.075 1.065 10.685 1.065 10.685 0.905 10.33 0.905 10.33 0.845 10.745 0.845 10.745 1.005 11.015 1.005 11.015 0.51 11.075 0.51 ;
      RECT 10.505 1.42 11.075 1.48 ;
      POLYGON 10.385 1.065 9.685 1.065 9.685 0.95 9.6 0.95 9.6 0.73 9.5 0.73 9.5 0.575 9.47 0.575 9.47 0.515 9.59 0.515 9.59 0.575 9.56 0.575 9.56 0.67 9.66 0.67 9.66 0.89 9.745 0.89 9.745 1.005 10.045 1.005 10.045 0.48 10.345 0.48 10.345 0.54 10.105 0.54 10.105 1.005 10.385 1.005 ;
      POLYGON 9.995 1.48 9.78 1.48 9.78 1.495 9.16 1.495 9.16 1.48 4.905 1.48 4.905 1.42 9.22 1.42 9.22 1.435 9.725 1.435 9.725 1.42 9.995 1.42 ;
      POLYGON 9.54 1.045 9.48 1.045 9.48 0.86 8.63 0.86 8.63 0.8 9.295 0.8 9.295 0.575 9.26 0.575 9.26 0.515 9.39 0.515 9.39 0.575 9.355 0.575 9.355 0.8 9.54 0.8 ;
      RECT 8.865 0.95 9.365 1.03 ;
      POLYGON 9.145 0.74 8.55 0.74 8.55 1.055 8.49 1.055 8.49 0.575 8.46 0.575 8.46 0.515 8.58 0.515 8.58 0.575 8.55 0.575 8.55 0.68 9.145 0.68 ;
      POLYGON 8.29 0.575 8.24 0.575 8.24 1.055 8.18 1.055 8.18 0.575 7.6 0.575 7.6 0.66 7.545 0.66 7.545 0.825 7.485 0.825 7.485 0.6 7.54 0.6 7.54 0.495 8.29 0.495 ;
      POLYGON 7.925 1.1 7.355 1.1 7.355 0.82 7.075 0.82 7.075 0.76 7.355 0.76 7.355 0.485 7.415 0.485 7.415 1.04 7.865 1.04 7.865 0.68 7.925 0.68 ;
      RECT 7.605 0.735 7.765 0.96 ;
      POLYGON 6.535 1.02 6.455 1.02 6.455 0.82 6.29 0.82 6.29 0.85 6.23 0.85 6.23 0.725 6.29 0.725 6.29 0.76 6.455 0.76 6.455 0.54 6.535 0.54 ;
      POLYGON 5.475 1.065 5.085 1.065 5.085 0.905 4.73 0.905 4.73 0.845 5.145 0.845 5.145 1.005 5.415 1.005 5.415 0.51 5.475 0.51 ;
      POLYGON 4.785 1.065 4.085 1.065 4.085 0.95 4 0.95 4 0.73 3.9 0.73 3.9 0.575 3.87 0.575 3.87 0.515 3.99 0.515 3.99 0.575 3.96 0.575 3.96 0.67 4.06 0.67 4.06 0.89 4.145 0.89 4.145 1.005 4.445 1.005 4.445 0.48 4.745 0.48 4.745 0.54 4.505 0.54 4.505 1.005 4.785 1.005 ;
      POLYGON 4.395 1.48 4.18 1.48 4.18 1.495 3.56 1.495 3.56 1.48 1.725 1.48 1.725 1.42 3.62 1.42 3.62 1.435 4.125 1.435 4.125 1.42 4.395 1.42 ;
      POLYGON 3.94 1.045 3.88 1.045 3.88 0.86 3.03 0.86 3.03 0.8 3.695 0.8 3.695 0.575 3.66 0.575 3.66 0.515 3.79 0.515 3.79 0.575 3.755 0.575 3.755 0.8 3.94 0.8 ;
      RECT 3.265 0.95 3.765 1.03 ;
      POLYGON 3.545 0.74 2.95 0.74 2.95 1.055 2.89 1.055 2.89 0.575 2.86 0.575 2.86 0.515 2.98 0.515 2.98 0.575 2.95 0.575 2.95 0.68 3.545 0.68 ;
      POLYGON 2.69 0.575 2.64 0.575 2.64 1.055 2.58 1.055 2.58 0.575 2 0.575 2 0.66 1.945 0.66 1.945 0.825 1.885 0.825 1.885 0.6 1.94 0.6 1.94 0.495 2.69 0.495 ;
      POLYGON 2.325 1.1 1.755 1.1 1.755 0.82 1.475 0.82 1.475 0.76 1.755 0.76 1.755 0.485 1.815 0.485 1.815 1.04 2.265 1.04 2.265 0.68 2.325 0.68 ;
      RECT 2.005 0.735 2.165 0.96 ;
      POLYGON 0.935 1.02 0.855 1.02 0.855 0.82 0.69 0.82 0.69 0.85 0.63 0.85 0.63 0.725 0.69 0.725 0.69 0.76 0.855 0.76 0.855 0.54 0.935 0.54 ;
  END
END SPDFF4RX2

MACRO SRDFFNQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SRDFFNQX1 0 0 ;
  SIZE 5.4 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 1.77 5.165 1.77 5.165 2.46 5.105 2.46 5.105 1.77 1.985 1.77 1.985 2.4 1.925 2.4 1.925 1.77 1.335 1.77 1.335 2.08 1.275 2.08 1.275 1.77 0 1.77 0 1.65 0.895 1.65 0.895 1.27 0.955 1.27 0.955 1.65 1.05 1.65 1.05 1.485 1.11 1.485 1.11 1.65 1.46 1.65 1.46 1.27 1.52 1.27 1.52 1.65 5.1 1.65 5.1 1.13 5.16 1.13 5.16 1.65 5.4 1.65 ;
    END
  END VDD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.065 2.585 2.06 2.585 2.06 2.605 1.825 2.605 1.825 2.465 2.06 2.465 2.06 2.525 2.065 2.525 ;
    END
  END SE
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.7 2.61 3.22 2.61 3.22 2 3.37 2 3.37 1.89 3.62 1.89 3.62 2 3.7 2 ;
    END
  END ExtVDD
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.579275 LAYER Metal1 ;
    ANTENNADIFFAREA 3.41475 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.22365 LAYER Metal1 ;
      ANTENNAMAXAREACAR 20.4751845 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 151.7102615 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.9 2.07 4.96 3.135 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.22 2.66 1.415 2.79 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 2.8 2.05 2.87 ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 3.48 0 3.48 0 3.36 0.855 3.36 0.855 2.97 0.915 2.97 0.915 3.36 1.305 3.36 1.305 2.94 1.365 2.94 1.365 3.36 1.925 3.36 1.925 2.96 1.985 2.96 1.985 3.36 3.22 3.36 3.22 3.025 3.28 3.025 3.28 3.36 3.64 3.36 3.64 3.025 3.7 3.025 3.7 3.36 5.105 3.36 5.105 2.875 5.165 2.875 5.165 3.36 5.4 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.4 0.06 5.16 0.06 5.16 0.465 5.1 0.465 5.1 0.06 3.755 0.06 3.755 0.57 3.695 0.57 3.695 0.06 1.315 0.06 1.315 0.465 1.255 0.465 1.255 0.06 0.955 0.06 0.955 0.465 0.895 0.465 0.895 0.06 0 0.06 0 -0.06 5.4 -0.06 ;
    END
  END VSS
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.775 2.52 0.985 2.645 ;
    END
  END CKN
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0441 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.361111 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 18.24074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.26 1.24 4.5 1.38 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 4.85 1.345 4.79 1.345 4.79 1.05 4.76 1.05 4.76 0.93 4.79 0.93 4.79 0.32 4.85 0.32 ;
      POLYGON 4.635 1.45 4.575 1.45 4.575 0.25 4.565 0.25 4.565 0.23 4.55 0.23 4.55 0.17 4.565 0.17 4.565 0.13 4.625 0.13 4.625 0.17 4.635 0.17 ;
      RECT 4.1 2.615 4.545 2.675 ;
      POLYGON 4.22 1.525 3.94 1.525 3.94 1.025 3.46 1.025 3.46 0.38 3.52 0.38 3.52 0.965 3.94 0.965 3.94 0.48 4 0.48 4 1.465 4.22 1.465 ;
      RECT 4.11 0.48 4.17 1.215 ;
      POLYGON 4.01 3.17 3.95 3.17 3.95 2.78 3.15 2.78 3.15 2.72 3.95 2.72 3.95 2 4.01 2 ;
      POLYGON 3.805 2.93 3.075 2.93 3.075 3.17 3.015 3.17 3.015 2 3.075 2 3.075 2.87 3.805 2.87 ;
      POLYGON 3.795 1.555 3.535 1.555 3.535 1.26 3.735 1.26 3.735 1.255 3.795 1.255 ;
      RECT 3.22 0.48 3.28 1.47 ;
      POLYGON 3.075 1.54 2.805 1.54 2.805 1.48 3.015 1.48 3.015 0.48 3.075 0.48 ;
      POLYGON 2.925 1.02 2.19 1.02 2.19 1.485 2.13 1.485 2.13 0.32 2.19 0.32 2.19 0.96 2.925 0.96 ;
      POLYGON 2.235 3.035 2.1 3.035 2.1 2.975 2.175 2.975 2.175 2.74 1.66 2.74 1.66 2.68 2.175 2.68 2.175 2.4 2.13 2.4 2.13 2.185 2.235 2.185 ;
      POLYGON 1.985 1.485 1.925 1.485 1.925 1.075 1.315 1.075 1.315 1.485 1.255 1.485 1.255 1.075 0.89 1.075 0.89 1.14 0.92 1.14 0.92 1.2 0.8 1.2 0.8 1.14 0.83 1.14 0.83 0.595 0.8 0.595 0.8 0.535 0.92 0.535 0.92 0.595 0.89 0.595 0.89 1.015 1.46 1.015 1.46 0.32 1.52 0.32 1.52 1.015 1.925 1.015 1.925 0.32 1.985 0.32 ;
      POLYGON 1.675 2.535 1.58 2.535 1.58 2.875 1.675 2.875 1.675 3.085 1.615 3.085 1.615 2.935 1.52 2.935 1.52 2.475 1.615 2.475 1.615 2.24 1.195 2.24 1.195 2.2 1.06 2.2 1.06 1.985 0.47 1.985 0.47 3.115 0.41 3.115 0.41 1.925 1.12 1.925 1.12 2.14 1.255 2.14 1.255 2.18 1.675 2.18 ;
      POLYGON 1.12 3.115 1.06 3.115 1.06 2.795 0.775 2.795 0.775 2.735 1.06 2.735 1.06 2.28 1.12 2.28 ;
      POLYGON 0.71 3.115 0.65 3.115 0.65 2.795 0.56 2.795 0.56 2.735 0.65 2.735 0.65 2.11 0.56 2.11 0.56 2.05 0.71 2.05 ;
      POLYGON 0.645 1.485 0.235 1.485 0.235 1.56 0.175 1.56 0.175 1.425 0.585 1.425 0.585 0.32 0.645 0.32 ;
      RECT 0.415 0.135 0.475 1.305 ;
      POLYGON 0.265 3.115 0.205 3.115 0.205 1.965 0.145 1.965 0.145 1.905 0.265 1.905 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END SRDFFNQX1

MACRO SRDFFNRQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SRDFFNRQX1 0 0 ;
  SIZE 5.6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 5.445 1.77 5.445 2.46 5.385 2.46 5.385 1.77 2.18 1.77 2.18 2.4 2.12 2.4 2.12 1.77 1.53 1.77 1.53 2.08 1.47 2.08 1.47 1.77 -0.005 1.77 -0.005 1.65 0.245 1.65 0.245 1.05 0.305 1.05 0.305 1.65 1.09 1.65 1.09 1.27 1.15 1.27 1.15 1.65 1.64 1.65 1.64 1.27 1.7 1.27 1.7 1.65 5.4 1.65 5.4 1.13 5.46 1.13 5.46 1.65 5.6 1.65 ;
    END
  END VDD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.26 2.585 2.255 2.585 2.255 2.605 2.02 2.605 2.02 2.465 2.255 2.465 2.255 2.525 2.26 2.525 ;
    END
  END SE
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.895 2.61 3.415 2.61 3.415 2 3.545 2 3.545 1.89 3.795 1.89 3.795 2 3.895 2 ;
    END
  END ExtVDD
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.5555555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.99 2.715 1.18 2.825 ;
    END
  END CKN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.385 0.905 0.375 0.905 0.375 0.98 0.245 0.98 0.245 0.74 0.375 0.74 0.375 0.845 0.385 0.845 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.955225 LAYER Metal1 ;
    ANTENNADIFFAREA 3.641925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.25605 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.35256775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 145.506737 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.24 3.135 5.18 3.135 5.18 2.86 5.01 2.86 5.01 2.655 5.18 2.655 5.18 2.07 5.24 2.07 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.9444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.415 2.66 1.61 2.84 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.97 2.8 2.225 2.88 ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 3.48 0 3.48 0 3.36 1.05 3.36 1.05 2.97 1.11 2.97 1.11 3.36 1.5 3.36 1.5 2.94 1.56 2.94 1.56 3.36 2.12 3.36 2.12 2.94 2.18 2.94 2.18 3.36 3.415 3.36 3.415 3.025 3.475 3.025 3.475 3.36 3.835 3.36 3.835 3.025 3.895 3.025 3.895 3.36 5.385 3.36 5.385 2.875 5.445 2.875 5.445 3.36 5.6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5.255 0.06 5.255 0.32 5.26 0.32 5.26 0.465 5.2 0.465 5.2 0.35 5.195 0.35 5.195 0.06 3.99 0.06 3.99 0.465 3.93 0.465 3.93 0.06 1.56 0.06 1.56 0.465 1.5 0.465 1.5 0.06 1.15 0.06 1.15 0.465 1.09 0.465 1.09 0.06 0.305 0.06 0.305 0.465 0.245 0.465 0.245 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.10185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.61 1.525 4.455 1.525 4.455 1.37 4.31 1.37 4.31 0.41 4.37 0.41 4.37 1.31 4.61 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.465 0.625 4.99 0.625 4.99 0.32 5.055 0.32 5.055 0.465 5.05 0.465 5.05 0.565 5.405 0.565 5.405 0.29 5.465 0.29 ;
      POLYGON 5.045 1.345 4.985 1.345 4.985 0.83 4.85 0.83 4.85 0.86 4.79 0.86 4.79 0.32 4.85 0.32 4.85 0.77 5.045 0.77 ;
      RECT 4.295 2.385 4.785 2.445 ;
      POLYGON 4.78 1.235 4.465 1.235 4.465 0.25 4.455 0.25 4.455 0.23 4.44 0.23 4.44 0.17 4.455 0.17 4.455 0.13 4.515 0.13 4.515 0.17 4.525 0.17 4.525 1.175 4.78 1.175 ;
      RECT 4.66 0.13 4.72 1.075 ;
      POLYGON 4.395 1.51 4.135 1.51 4.135 0.83 3.6 0.83 3.6 0.245 3.66 0.245 3.66 0.77 4.135 0.77 4.135 0.32 4.195 0.32 4.195 1.45 4.395 1.45 ;
      POLYGON 4.205 3.17 4.145 3.17 4.145 2.78 3.345 2.78 3.345 2.72 4.145 2.72 4.145 2 4.205 2 ;
      POLYGON 4 2.93 3.27 2.93 3.27 3.17 3.21 3.17 3.21 2 3.27 2 3.27 2.87 4 2.87 ;
      RECT 3.71 1.24 3.99 1.525 ;
      RECT 3.415 0.32 3.475 1.455 ;
      POLYGON 3.27 1.52 2.935 1.52 2.935 1.46 3.21 1.46 3.21 0.32 3.27 0.32 ;
      RECT 2.675 0.6 2.735 1.29 ;
      POLYGON 2.445 0.83 2.385 0.83 2.385 1.485 2.325 1.485 2.325 0.32 2.385 0.32 2.385 0.77 2.445 0.77 ;
      POLYGON 2.385 3.085 2.325 3.085 2.325 2.74 1.855 2.74 1.855 2.68 2.325 2.68 2.325 2.185 2.385 2.185 ;
      POLYGON 2.18 1.485 2.12 1.485 2.12 0.585 1.39 0.585 1.39 1.485 1.33 1.485 1.33 0.585 1.115 0.585 1.115 0.595 1.085 0.595 1.085 1.14 1.115 1.14 1.115 1.2 0.995 1.2 0.995 1.14 1.025 1.14 1.025 0.595 0.995 0.595 0.995 0.535 1.025 0.535 1.025 0.525 1.295 0.525 1.295 0.32 1.355 0.32 1.355 0.525 2.12 0.525 2.12 0.32 2.18 0.32 ;
      POLYGON 1.87 2.535 1.745 2.535 1.745 2.875 1.87 2.875 1.87 3.085 1.81 3.085 1.81 2.935 1.685 2.935 1.685 2.475 1.81 2.475 1.81 2.24 1.39 2.24 1.39 2.2 1.255 2.2 1.255 1.985 0.665 1.985 0.665 3.115 0.605 3.115 0.605 1.925 1.315 1.925 1.315 2.14 1.45 2.14 1.45 2.18 1.87 2.18 ;
      POLYGON 1.315 3.115 1.255 3.115 1.255 2.64 0.945 2.64 0.945 2.58 1.255 2.58 1.255 2.28 1.315 2.28 ;
      POLYGON 0.905 2.51 0.795 2.51 0.795 2.97 0.905 2.97 0.905 3.115 0.845 3.115 0.845 3.03 0.735 3.03 0.735 2.45 0.845 2.45 0.845 2.105 0.77 2.105 0.77 2.045 0.905 2.045 ;
      POLYGON 0.84 1.485 0.43 1.485 0.43 1.56 0.37 1.56 0.37 1.425 0.78 1.425 0.78 0.32 0.84 0.32 ;
      RECT 0.61 0.135 0.67 1.305 ;
      POLYGON 0.55 0.985 0.51 0.985 0.51 1.265 0.45 1.265 0.45 0.32 0.51 0.32 0.51 0.865 0.55 0.865 ;
      POLYGON 0.46 3.115 0.4 3.115 0.4 1.965 0.34 1.965 0.34 1.905 0.46 1.905 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END SRDFFNRQX1

MACRO SRDFFNRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SRDFFNRX1 0 0 ;
  SIZE 6.2 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 5.93 1.77 5.93 2.46 5.87 2.46 5.87 1.77 5.25 1.77 5.25 2.48 5.19 2.48 5.19 1.77 2.18 1.77 2.18 2.4 2.12 2.4 2.12 1.77 1.53 1.77 1.53 2.08 1.47 2.08 1.47 1.77 0 1.77 0 1.65 0.245 1.65 0.245 1.05 0.305 1.05 0.305 1.65 1.09 1.65 1.09 1.27 1.15 1.27 1.15 1.65 1.745 1.65 1.745 1.27 1.805 1.27 1.805 1.65 5.43 1.65 5.43 1.13 5.49 1.13 5.49 1.65 6.2 1.65 ;
    END
  END VDD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.26 2.585 2.255 2.585 2.255 2.605 2.02 2.605 2.02 2.465 2.255 2.465 2.255 2.525 2.26 2.525 ;
    END
  END SE
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.895 2.61 3.415 2.61 3.415 2 3.545 2 3.545 1.89 3.795 1.89 3.795 2 3.895 2 ;
    END
  END ExtVDD
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.5555555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.99 2.715 1.18 2.825 ;
    END
  END CKN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.385 0.905 0.375 0.905 0.375 0.98 0.245 0.98 0.245 0.74 0.375 0.74 0.375 0.845 0.385 0.845 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4337 LAYER Metal1 ;
    ANTENNADIFFAREA 4.111775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3015 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.02222225 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 135.83084575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.77 2.84 5.725 2.84 5.725 3.135 5.665 3.135 5.665 2.84 5.605 2.84 5.605 2.66 5.665 2.66 5.665 2.07 5.725 2.07 5.725 2.66 5.77 2.66 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4337 LAYER Metal1 ;
    ANTENNADIFFAREA 4.111775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3015 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.02222225 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 135.83084575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.045 3.13 4.985 3.13 4.985 2.85 4.805 2.85 4.805 2.655 4.985 2.655 4.985 2.09 5.045 2.09 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.9444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.415 2.66 1.61 2.84 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.97 2.8 2.225 2.88 ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 3.48 0 3.48 0 3.36 1.05 3.36 1.05 2.97 1.11 2.97 1.11 3.36 1.5 3.36 1.5 2.94 1.56 2.94 1.56 3.36 2.12 3.36 2.12 2.94 2.18 2.94 2.18 3.36 3.415 3.36 3.415 3.025 3.475 3.025 3.475 3.36 3.835 3.36 3.835 3.025 3.895 3.025 3.895 3.36 5.19 3.36 5.19 2.87 5.25 2.87 5.25 3.36 5.87 3.36 5.87 2.875 5.93 2.875 5.93 3.36 6.2 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 5.86 0.06 5.86 0.465 5.8 0.465 5.8 0.06 5.45 0.06 5.45 0.465 5.39 0.465 5.39 0.06 3.99 0.06 3.99 0.465 3.93 0.465 3.93 0.06 1.84 0.06 1.84 0.465 1.78 0.465 1.78 0.06 1.15 0.06 1.15 0.465 1.09 0.465 1.09 0.06 0.305 0.06 0.305 0.465 0.245 0.465 0.245 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.10185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.61 1.525 4.455 1.525 4.455 1.37 4.31 1.37 4.31 0.41 4.37 0.41 4.37 1.31 4.61 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.8 1.345 5.74 1.345 5.74 1.015 5.25 1.015 5.25 1.345 5.19 1.345 5.19 0.955 5.8 0.955 ;
      POLYGON 5.655 0.67 5.19 0.67 5.19 0.32 5.25 0.32 5.25 0.61 5.595 0.61 5.595 0.32 5.655 0.32 ;
      POLYGON 5.485 3.07 5.425 3.07 5.425 2.71 5.13 2.71 5.13 2.65 5.425 2.65 5.425 2.175 5.485 2.175 ;
      RECT 4.985 0.32 5.045 1.345 ;
      POLYGON 4.81 1.07 4.465 1.07 4.465 0.25 4.455 0.25 4.455 0.23 4.44 0.23 4.44 0.17 4.455 0.17 4.455 0.13 4.515 0.13 4.515 0.17 4.525 0.17 4.525 1.01 4.81 1.01 ;
      RECT 4.295 2.385 4.74 2.445 ;
      POLYGON 4.395 1.51 4.135 1.51 4.135 0.83 3.6 0.83 3.6 0.245 3.66 0.245 3.66 0.77 4.135 0.77 4.135 0.32 4.195 0.32 4.195 1.45 4.395 1.45 ;
      POLYGON 4.205 3.17 4.145 3.17 4.145 2.78 3.345 2.78 3.345 2.72 4.145 2.72 4.145 2 4.205 2 ;
      POLYGON 4 2.93 3.27 2.93 3.27 3.17 3.21 3.17 3.21 2 3.27 2 3.27 2.87 4 2.87 ;
      RECT 3.71 1.24 3.99 1.525 ;
      RECT 3.415 0.32 3.475 1.455 ;
      POLYGON 3.27 1.52 2.935 1.52 2.935 1.46 3.21 1.46 3.21 0.32 3.27 0.32 ;
      RECT 2.675 0.6 2.735 1.29 ;
      POLYGON 2.385 3.085 2.325 3.085 2.325 2.74 1.855 2.74 1.855 2.68 2.325 2.68 2.325 2.185 2.385 2.185 ;
      POLYGON 2.31 0.83 2.25 0.83 2.25 1.485 2.19 1.485 2.19 0.32 2.25 0.32 2.25 0.77 2.31 0.77 ;
      POLYGON 2.045 1.485 1.985 1.485 1.985 0.585 1.495 0.585 1.495 1.485 1.435 1.485 1.435 0.585 1.115 0.585 1.115 0.595 1.085 0.595 1.085 1.14 1.115 1.14 1.115 1.2 0.995 1.2 0.995 1.14 1.025 1.14 1.025 0.595 0.995 0.595 0.995 0.535 1.025 0.535 1.025 0.525 1.295 0.525 1.295 0.32 1.355 0.32 1.355 0.525 1.985 0.525 1.985 0.32 2.045 0.32 ;
      POLYGON 1.87 2.535 1.745 2.535 1.745 2.875 1.87 2.875 1.87 3.085 1.81 3.085 1.81 2.935 1.685 2.935 1.685 2.475 1.81 2.475 1.81 2.24 1.39 2.24 1.39 2.2 1.255 2.2 1.255 1.985 0.665 1.985 0.665 3.115 0.605 3.115 0.605 1.925 1.315 1.925 1.315 2.14 1.45 2.14 1.45 2.18 1.87 2.18 ;
      POLYGON 1.315 3.115 1.255 3.115 1.255 2.64 0.945 2.64 0.945 2.58 1.255 2.58 1.255 2.28 1.315 2.28 ;
      RECT 1.19 0.68 1.25 1.09 ;
      POLYGON 0.905 2.51 0.795 2.51 0.795 2.97 0.905 2.97 0.905 3.115 0.845 3.115 0.845 3.03 0.735 3.03 0.735 2.45 0.845 2.45 0.845 2.105 0.77 2.105 0.77 2.045 0.905 2.045 ;
      POLYGON 0.84 1.485 0.43 1.485 0.43 1.56 0.37 1.56 0.37 1.425 0.78 1.425 0.78 0.32 0.84 0.32 ;
      RECT 0.61 0.135 0.67 1.305 ;
      POLYGON 0.55 0.95 0.51 0.95 0.51 1.265 0.45 1.265 0.45 0.32 0.51 0.32 0.51 0.83 0.55 0.83 ;
      POLYGON 0.46 3.115 0.4 3.115 0.4 1.965 0.34 1.965 0.34 1.905 0.46 1.905 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END SRDFFNRX1

MACRO SRDFFNSQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SRDFFNSQX1 0 0 ;
  SIZE 6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 1.77 5.625 1.77 5.625 2.46 5.565 2.46 5.565 1.77 1.98 1.77 1.98 2.4 1.92 2.4 1.92 1.77 1.33 1.77 1.33 2.08 1.27 2.08 1.27 1.77 -0.005 1.77 -0.005 1.65 0.89 1.65 0.89 1.27 0.95 1.27 0.95 1.65 1.045 1.65 1.045 1.27 1.105 1.27 1.105 1.65 1.455 1.65 1.455 1.27 1.515 1.27 1.515 1.65 5.23 1.65 5.23 1.13 5.29 1.13 5.29 1.65 5.64 1.65 5.64 1.13 5.7 1.13 5.7 1.65 6 1.65 ;
    END
  END VDD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.14814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.06 2.585 2.055 2.585 2.055 2.605 1.82 2.605 1.82 2.505 2.055 2.505 2.055 2.525 2.06 2.525 ;
    END
  END SE
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0516 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.5925925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 23.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.165 0.96 1.105 0.96 1.105 1.14 1.135 1.14 1.135 1.2 1.015 1.2 1.015 1.14 1.045 1.14 1.045 0.96 1.025 0.96 1.025 0.72 1.165 0.72 ;
    END
  END SN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.695 2.61 3.215 2.61 3.215 2 3.345 2 3.345 1.89 3.595 1.89 3.595 2 3.695 2 ;
    END
  END ExtVDD
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.64814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.805 2.715 0.98 2.845 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.983575 LAYER Metal1 ;
    ANTENNADIFFAREA 3.716825 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.22365 LAYER Metal1 ;
      ANTENNAMAXAREACAR 22.28291975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 164.06438625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.42 3.135 5.36 3.135 5.36 2.855 5.21 2.855 5.21 2.65 5.36 2.65 5.36 2.07 5.42 2.07 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.85185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 2.66 1.41 2.835 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.77 2.8 2.025 2.88 ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 3.48 0 3.48 0 3.36 0.85 3.36 0.85 2.97 0.91 2.97 0.91 3.36 1.3 3.36 1.3 2.94 1.36 2.94 1.36 3.36 1.92 3.36 1.92 2.94 1.98 2.94 1.98 3.36 3.215 3.36 3.215 3.025 3.275 3.025 3.275 3.36 3.635 3.36 3.635 3.025 3.695 3.025 3.695 3.36 5.565 3.36 5.565 2.875 5.625 2.875 5.625 3.36 6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6 0.06 5.265 0.06 5.265 0.35 5.26 0.35 5.26 0.465 5.2 0.465 5.2 0.32 5.205 0.32 5.205 0.06 3.79 0.06 3.79 0.465 3.73 0.465 3.73 0.06 0.95 0.06 0.95 0.32 1.125 0.32 1.125 0.465 0.89 0.465 0.89 0.06 0 0.06 0 -0.06 6 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.10185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.41 1.525 4.255 1.525 4.255 1.37 4.11 1.37 4.11 0.41 4.17 0.41 4.17 1.31 4.41 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.495 1.345 5.435 1.345 5.435 1.015 5.05 1.015 5.05 1.345 4.99 1.345 4.99 0.955 5.495 0.955 ;
      RECT 4.785 0.32 4.845 1.345 ;
      RECT 4.095 2.385 4.54 2.445 ;
      POLYGON 4.535 1.13 4.265 1.13 4.265 0.25 4.255 0.25 4.255 0.23 4.24 0.23 4.24 0.17 4.255 0.17 4.255 0.13 4.315 0.13 4.315 0.17 4.325 0.17 4.325 1.07 4.535 1.07 ;
      RECT 4.445 0.135 4.505 0.995 ;
      POLYGON 4.195 1.51 3.935 1.51 3.935 0.83 3.4 0.83 3.4 0.245 3.46 0.245 3.46 0.77 3.935 0.77 3.935 0.32 3.995 0.32 3.995 1.45 4.195 1.45 ;
      POLYGON 4.005 3.17 3.945 3.17 3.945 2.78 3.145 2.78 3.145 2.72 3.945 2.72 3.945 2 4.005 2 ;
      POLYGON 3.8 2.93 3.07 2.93 3.07 3.17 3.01 3.17 3.01 2 3.07 2 3.07 2.87 3.8 2.87 ;
      RECT 3.51 1.24 3.79 1.525 ;
      RECT 3.215 0.32 3.275 1.455 ;
      POLYGON 3.07 1.52 2.735 1.52 2.735 1.46 3.01 1.46 3.01 0.32 3.07 0.32 ;
      RECT 2.475 0.6 2.535 1.29 ;
      POLYGON 2.245 0.83 2.185 0.83 2.185 1.485 2.125 1.485 2.125 0.32 2.185 0.32 2.185 0.77 2.245 0.77 ;
      POLYGON 2.185 3.085 2.125 3.085 2.125 2.74 1.655 2.74 1.655 2.68 2.125 2.68 2.125 2.185 2.185 2.185 ;
      POLYGON 1.98 1.485 1.92 1.485 1.92 0.585 1.31 0.585 1.31 1.485 1.25 1.485 1.25 0.585 0.915 0.585 0.915 0.595 0.885 0.595 0.885 1.14 0.915 1.14 0.915 1.2 0.795 1.2 0.795 1.14 0.825 1.14 0.825 0.595 0.795 0.595 0.795 0.535 0.825 0.535 0.825 0.525 1.375 0.525 1.375 0.32 1.435 0.32 1.435 0.525 1.92 0.525 1.92 0.32 1.98 0.32 ;
      POLYGON 1.67 2.535 1.545 2.535 1.545 2.875 1.67 2.875 1.67 3.085 1.61 3.085 1.61 2.935 1.485 2.935 1.485 2.475 1.61 2.475 1.61 2.21 1.145 2.21 1.145 2.18 1.055 2.18 1.055 1.985 0.465 1.985 0.465 3.115 0.405 3.115 0.405 1.925 1.115 1.925 1.115 2.12 1.205 2.12 1.205 2.15 1.67 2.15 ;
      RECT 1.38 0.67 1.44 1.13 ;
      POLYGON 1.115 3.115 1.055 3.115 1.055 2.64 0.745 2.64 0.745 2.58 1.055 2.58 1.055 2.28 1.115 2.28 ;
      POLYGON 0.705 2.51 0.595 2.51 0.595 2.97 0.705 2.97 0.705 3.115 0.645 3.115 0.645 3.03 0.535 3.03 0.535 2.45 0.645 2.45 0.645 2.105 0.57 2.105 0.57 2.045 0.705 2.045 ;
      POLYGON 0.64 1.485 0.23 1.485 0.23 1.56 0.17 1.56 0.17 1.425 0.58 1.425 0.58 0.32 0.64 0.32 ;
      RECT 0.41 0.135 0.47 1.305 ;
      POLYGON 0.26 3.115 0.2 3.115 0.2 1.965 0.14 1.965 0.14 1.905 0.26 1.905 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END SRDFFNSQX1

MACRO SRDFFNSRQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SRDFFNSRQX1 0 0 ;
  SIZE 6.2 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 5.93 1.77 5.93 2.46 5.87 2.46 5.87 1.77 2.18 1.77 2.18 2.4 2.12 2.4 2.12 1.77 1.53 1.77 1.53 2.08 1.47 2.08 1.47 1.77 -0.005 1.77 -0.005 1.65 0.245 1.65 0.245 1.05 0.305 1.05 0.305 1.65 1.09 1.65 1.09 1.27 1.15 1.27 1.15 1.65 1.88 1.65 1.88 1.27 1.94 1.27 1.94 1.65 5.43 1.65 5.43 1.13 5.49 1.13 5.49 1.65 5.945 1.65 5.945 1.13 6.005 1.13 6.005 1.65 6.2 1.65 ;
    END
  END VDD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.26 2.585 2.255 2.585 2.255 2.605 2.02 2.605 2.02 2.465 2.255 2.465 2.255 2.525 2.26 2.525 ;
    END
  END SE
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0516 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.5925925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 23.37962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.355 0.84 1.29 0.84 1.29 1.14 1.32 1.14 1.32 1.2 1.2 1.2 1.2 1.14 1.23 1.14 1.23 0.84 1.21 0.84 1.21 0.72 1.355 0.72 ;
    END
  END SN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.895 2.61 3.415 2.61 3.415 2 3.545 2 3.545 1.89 3.795 1.89 3.795 2 3.895 2 ;
    END
  END ExtVDD
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.22222225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.18 2.825 0.9 2.825 0.9 2.715 1.16 2.715 1.16 2.765 1.18 2.765 ;
    END
  END CKN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.66666675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.385 0.905 0.375 0.905 0.375 0.98 0.265 0.98 0.265 0.74 0.375 0.74 0.375 0.845 0.385 0.845 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.429625 LAYER Metal1 ;
    ANTENNADIFFAREA 3.9912 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.25605 LAYER Metal1 ;
      ANTENNAMAXAREACAR 21.205331 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 159.062683 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.665 2.07 5.725 3.135 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.415 2.66 1.61 2.79 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.95 2.8 2.245 2.87 ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 3.48 0 3.48 0 3.36 1.05 3.36 1.05 2.97 1.11 2.97 1.11 3.36 1.5 3.36 1.5 2.94 1.56 2.94 1.56 3.36 2.12 3.36 2.12 2.94 2.18 2.94 2.18 3.36 3.415 3.36 3.415 3.025 3.475 3.025 3.475 3.36 3.835 3.36 3.835 3.025 3.895 3.025 3.895 3.36 5.87 3.36 5.87 2.875 5.93 2.875 5.93 3.36 6.2 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 6.065 0.06 6.065 0.465 6.005 0.465 6.005 0.06 3.99 0.06 3.99 0.465 3.93 0.465 3.93 0.06 1.15 0.06 1.15 0.32 1.325 0.32 1.325 0.465 1.09 0.465 1.09 0.06 0.305 0.06 0.305 0.465 0.245 0.465 0.245 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.10185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.61 1.525 4.455 1.525 4.455 1.37 4.31 1.37 4.31 0.41 4.37 0.41 4.37 1.31 4.61 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.86 0.465 5.8 0.465 5.8 0.26 5.45 0.26 5.45 0.465 5.39 0.465 5.39 0.2 5.86 0.2 ;
      POLYGON 5.8 1.345 5.74 1.345 5.74 1.015 5.25 1.015 5.25 1.345 5.19 1.345 5.19 0.955 5.8 0.955 ;
      POLYGON 5.655 0.67 5.19 0.67 5.19 0.32 5.25 0.32 5.25 0.61 5.595 0.61 5.595 0.32 5.655 0.32 ;
      RECT 4.985 0.32 5.045 1.345 ;
      RECT 4.295 2.385 4.74 2.445 ;
      POLYGON 4.735 1.13 4.465 1.13 4.465 0.25 4.455 0.25 4.455 0.23 4.44 0.23 4.44 0.17 4.455 0.17 4.455 0.13 4.515 0.13 4.515 0.17 4.525 0.17 4.525 1.07 4.735 1.07 ;
      RECT 4.645 0.135 4.705 0.995 ;
      POLYGON 4.395 1.51 4.135 1.51 4.135 0.83 3.6 0.83 3.6 0.245 3.66 0.245 3.66 0.77 4.135 0.77 4.135 0.32 4.195 0.32 4.195 1.45 4.395 1.45 ;
      POLYGON 4.205 3.17 4.145 3.17 4.145 2.78 3.345 2.78 3.345 2.72 4.145 2.72 4.145 2 4.205 2 ;
      POLYGON 4 2.93 3.27 2.93 3.27 3.17 3.21 3.17 3.21 2 3.27 2 3.27 2.87 4 2.87 ;
      RECT 3.71 1.24 3.99 1.525 ;
      RECT 3.415 0.32 3.475 1.455 ;
      POLYGON 3.27 1.52 2.935 1.52 2.935 1.46 3.21 1.46 3.21 0.32 3.27 0.32 ;
      RECT 2.675 0.6 2.735 1.29 ;
      POLYGON 2.445 0.83 2.385 0.83 2.385 1.485 2.325 1.485 2.325 0.32 2.385 0.32 2.385 0.77 2.445 0.77 ;
      POLYGON 2.385 3.085 2.325 3.085 2.325 2.74 1.855 2.74 1.855 2.68 2.325 2.68 2.325 2.185 2.385 2.185 ;
      POLYGON 2.265 1.19 2.18 1.19 2.18 1.485 2.12 1.485 2.12 1.13 2.205 1.13 2.205 0.585 1.51 0.585 1.51 1.27 1.63 1.27 1.63 1.485 1.295 1.485 1.295 1.27 1.45 1.27 1.45 0.585 1.115 0.585 1.115 0.595 1.085 0.595 1.085 1.14 1.115 1.14 1.115 1.2 0.995 1.2 0.995 1.14 1.025 1.14 1.025 0.595 0.995 0.595 0.995 0.535 1.025 0.535 1.025 0.525 1.675 0.525 1.675 0.32 1.735 0.32 1.735 0.525 2.12 0.525 2.12 0.32 2.18 0.32 2.18 0.525 2.265 0.525 ;
      POLYGON 2.115 0.705 2.075 0.705 2.075 0.75 2.06 0.75 2.06 1.18 2 1.18 2 0.705 1.995 0.705 1.995 0.645 2.115 0.645 ;
      POLYGON 1.975 0.465 1.915 0.465 1.915 0.255 1.53 0.255 1.53 0.465 1.47 0.465 1.47 0.195 1.975 0.195 ;
      POLYGON 1.915 0.705 1.885 0.705 1.885 1.185 1.725 1.185 1.725 1.2 1.605 1.2 1.605 1.14 1.635 1.14 1.635 1.125 1.825 1.125 1.825 0.705 1.795 0.705 1.795 0.645 1.915 0.645 ;
      POLYGON 1.87 2.535 1.745 2.535 1.745 2.875 1.87 2.875 1.87 3.085 1.81 3.085 1.81 2.935 1.685 2.935 1.685 2.475 1.81 2.475 1.81 2.24 1.39 2.24 1.39 2.2 1.255 2.2 1.255 1.985 0.665 1.985 0.665 3.115 0.605 3.115 0.605 1.925 1.315 1.925 1.315 2.14 1.45 2.14 1.45 2.18 1.87 2.18 ;
      POLYGON 1.315 3.115 1.255 3.115 1.255 2.64 0.945 2.64 0.945 2.58 1.255 2.58 1.255 2.28 1.315 2.28 ;
      POLYGON 0.905 2.51 0.795 2.51 0.795 2.97 0.905 2.97 0.905 3.115 0.845 3.115 0.845 3.03 0.735 3.03 0.735 2.45 0.845 2.45 0.845 2.105 0.77 2.105 0.77 2.045 0.905 2.045 ;
      POLYGON 0.84 1.485 0.43 1.485 0.43 1.56 0.37 1.56 0.37 1.425 0.78 1.425 0.78 0.32 0.84 0.32 ;
      RECT 0.61 0.135 0.67 1.305 ;
      POLYGON 0.55 0.985 0.51 0.985 0.51 1.265 0.45 1.265 0.45 0.32 0.51 0.32 0.51 0.865 0.55 0.865 ;
      POLYGON 0.46 3.115 0.4 3.115 0.4 1.965 0.34 1.965 0.34 1.905 0.46 1.905 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END SRDFFNSRQX1

MACRO SRDFFNSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SRDFFNSRX1 0 0 ;
  SIZE 6.2 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 5.93 1.77 5.93 2.46 5.87 2.46 5.87 1.77 5.25 1.77 5.25 2.48 5.19 2.48 5.19 1.77 2.18 1.77 2.18 2.4 2.12 2.4 2.12 1.77 1.53 1.77 1.53 2.08 1.47 2.08 1.47 1.77 -0.005 1.77 -0.005 1.65 0.245 1.65 0.245 1.05 0.305 1.05 0.305 1.65 1.09 1.65 1.09 1.27 1.15 1.27 1.15 1.65 1.88 1.65 1.88 1.27 1.94 1.27 1.94 1.65 5.43 1.65 5.43 1.13 5.49 1.13 5.49 1.65 5.945 1.65 5.945 1.13 6.005 1.13 6.005 1.65 6.2 1.65 ;
    END
  END VDD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.24074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.035 2.48 2.26 2.605 ;
    END
  END SE
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1045 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 3.22530875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 30 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.37 0.925 1.29 0.925 1.29 1.14 1.32 1.14 1.32 1.2 1.2 1.2 1.2 1.14 1.23 1.14 1.23 0.925 1.21 0.925 1.21 0.72 1.37 0.72 ;
    END
  END SN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.895 2.61 3.415 2.61 3.415 2 3.545 2 3.545 1.89 3.795 1.89 3.795 2 3.895 2 ;
    END
  END ExtVDD
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.01 2.69 1.18 2.845 ;
    END
  END CKN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.4814815 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.385 0.905 0.375 0.905 0.375 0.95 0.245 0.95 0.245 0.74 0.375 0.74 0.375 0.845 0.385 0.845 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.683475 LAYER Metal1 ;
    ANTENNADIFFAREA 4.2416 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3015 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.85066325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 142.60696525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.765 2.835 5.725 2.835 5.725 3.135 5.665 3.135 5.665 2.835 5.635 2.835 5.635 2.48 5.665 2.48 5.665 2.07 5.725 2.07 5.725 2.48 5.765 2.48 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.683475 LAYER Metal1 ;
    ANTENNADIFFAREA 4.271325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3015 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.85066325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 142.60696525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.045 3.13 4.985 3.13 4.985 2.825 4.825 2.825 4.825 2.68 4.985 2.68 4.985 2.09 5.045 2.09 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.415 2.68 1.61 2.82 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.97 2.8 2.225 2.88 ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 3.48 0 3.48 0 3.36 1.05 3.36 1.05 2.97 1.11 2.97 1.11 3.36 1.5 3.36 1.5 2.94 1.56 2.94 1.56 3.36 2.12 3.36 2.12 2.94 2.18 2.94 2.18 3.36 3.415 3.36 3.415 3.025 3.475 3.025 3.475 3.36 3.835 3.36 3.835 3.025 3.895 3.025 3.895 3.36 5.19 3.36 5.19 2.87 5.25 2.87 5.25 3.36 5.87 3.36 5.87 2.875 5.93 2.875 5.93 3.36 6.2 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 6.065 0.06 6.065 0.465 6.005 0.465 6.005 0.06 3.99 0.06 3.99 0.465 3.93 0.465 3.93 0.06 1.15 0.06 1.15 0.32 1.325 0.32 1.325 0.465 1.09 0.465 1.09 0.06 0.305 0.06 0.305 0.465 0.245 0.465 0.245 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.10185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.61 1.525 4.455 1.525 4.455 1.37 4.31 1.37 4.31 0.41 4.37 0.41 4.37 1.31 4.61 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.86 0.465 5.8 0.465 5.8 0.26 5.45 0.26 5.45 0.465 5.39 0.465 5.39 0.2 5.86 0.2 ;
      POLYGON 5.8 1.345 5.74 1.345 5.74 1.015 5.25 1.015 5.25 1.345 5.19 1.345 5.19 0.955 5.8 0.955 ;
      POLYGON 5.655 0.67 5.19 0.67 5.19 0.32 5.25 0.32 5.25 0.61 5.595 0.61 5.595 0.32 5.655 0.32 ;
      POLYGON 5.485 3.07 5.425 3.07 5.425 2.71 5.13 2.71 5.13 2.65 5.425 2.65 5.425 2.175 5.485 2.175 ;
      RECT 4.985 0.32 5.045 1.345 ;
      RECT 4.295 2.385 4.74 2.445 ;
      POLYGON 4.735 1.13 4.465 1.13 4.465 0.25 4.455 0.25 4.455 0.23 4.44 0.23 4.44 0.17 4.455 0.17 4.455 0.13 4.515 0.13 4.515 0.17 4.525 0.17 4.525 1.07 4.735 1.07 ;
      RECT 4.645 0.135 4.705 0.995 ;
      POLYGON 4.395 1.51 4.135 1.51 4.135 0.83 3.6 0.83 3.6 0.245 3.66 0.245 3.66 0.77 4.135 0.77 4.135 0.32 4.195 0.32 4.195 1.45 4.395 1.45 ;
      POLYGON 4.205 3.17 4.145 3.17 4.145 2.78 3.345 2.78 3.345 2.72 4.145 2.72 4.145 2 4.205 2 ;
      POLYGON 4 2.93 3.27 2.93 3.27 3.17 3.21 3.17 3.21 2 3.27 2 3.27 2.87 4 2.87 ;
      RECT 3.71 1.24 3.99 1.525 ;
      RECT 3.415 0.32 3.475 1.455 ;
      POLYGON 3.27 1.52 2.935 1.52 2.935 1.46 3.21 1.46 3.21 0.32 3.27 0.32 ;
      RECT 2.675 0.6 2.735 1.29 ;
      POLYGON 2.445 0.83 2.385 0.83 2.385 1.485 2.325 1.485 2.325 0.32 2.385 0.32 2.385 0.77 2.445 0.77 ;
      POLYGON 2.385 3.085 2.325 3.085 2.325 2.74 1.855 2.74 1.855 2.68 2.325 2.68 2.325 2.185 2.385 2.185 ;
      POLYGON 2.265 1.19 2.18 1.19 2.18 1.485 2.12 1.485 2.12 1.13 2.205 1.13 2.205 0.585 1.51 0.585 1.51 1.27 1.63 1.27 1.63 1.485 1.295 1.485 1.295 1.27 1.45 1.27 1.45 0.585 1.115 0.585 1.115 0.595 1.085 0.595 1.085 1.14 1.115 1.14 1.115 1.2 0.995 1.2 0.995 1.14 1.025 1.14 1.025 0.595 0.995 0.595 0.995 0.535 1.025 0.535 1.025 0.525 1.675 0.525 1.675 0.32 1.735 0.32 1.735 0.525 2.12 0.525 2.12 0.32 2.18 0.32 2.18 0.525 2.265 0.525 ;
      POLYGON 2.115 0.705 2.075 0.705 2.075 0.75 2.06 0.75 2.06 1.18 2 1.18 2 0.705 1.995 0.705 1.995 0.645 2.115 0.645 ;
      POLYGON 1.975 0.465 1.915 0.465 1.915 0.255 1.53 0.255 1.53 0.465 1.47 0.465 1.47 0.195 1.975 0.195 ;
      POLYGON 1.915 0.705 1.885 0.705 1.885 1.185 1.725 1.185 1.725 1.2 1.605 1.2 1.605 1.14 1.635 1.14 1.635 1.125 1.825 1.125 1.825 0.705 1.795 0.705 1.795 0.645 1.915 0.645 ;
      POLYGON 1.87 2.535 1.745 2.535 1.745 2.875 1.87 2.875 1.87 3.085 1.81 3.085 1.81 2.935 1.685 2.935 1.685 2.475 1.81 2.475 1.81 2.24 1.39 2.24 1.39 2.2 1.255 2.2 1.255 1.985 0.665 1.985 0.665 3.115 0.605 3.115 0.605 1.925 1.315 1.925 1.315 2.14 1.45 2.14 1.45 2.18 1.87 2.18 ;
      POLYGON 1.315 3.115 1.255 3.115 1.255 2.61 0.945 2.61 0.945 2.55 1.255 2.55 1.255 2.28 1.315 2.28 ;
      POLYGON 0.905 2.49 0.795 2.49 0.795 2.97 0.905 2.97 0.905 3.115 0.845 3.115 0.845 3.03 0.735 3.03 0.735 2.43 0.845 2.43 0.845 2.105 0.77 2.105 0.77 2.045 0.905 2.045 ;
      POLYGON 0.84 1.485 0.43 1.485 0.43 1.56 0.37 1.56 0.37 1.425 0.78 1.425 0.78 0.32 0.84 0.32 ;
      RECT 0.61 0.135 0.67 1.305 ;
      POLYGON 0.55 0.985 0.51 0.985 0.51 1.265 0.45 1.265 0.45 0.32 0.51 0.32 0.51 0.865 0.55 0.865 ;
      POLYGON 0.46 3.115 0.4 3.115 0.4 1.965 0.34 1.965 0.34 1.905 0.46 1.905 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END SRDFFNSRX1

MACRO SRDFFNSX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SRDFFNSX1 0 0 ;
  SIZE 6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 1.77 5.73 1.77 5.73 2.46 5.67 2.46 5.67 1.77 5.05 1.77 5.05 2.48 4.99 2.48 4.99 1.77 1.98 1.77 1.98 2.4 1.92 2.4 1.92 1.77 1.33 1.77 1.33 2.08 1.27 2.08 1.27 1.77 -0.005 1.77 -0.005 1.65 0.89 1.65 0.89 1.27 0.95 1.27 0.95 1.65 1.575 1.65 1.575 1.27 1.635 1.27 1.635 1.65 5.23 1.65 5.23 1.13 5.29 1.13 5.29 1.65 5.64 1.65 5.64 1.13 5.7 1.13 5.7 1.65 6 1.65 ;
    END
  END VDD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.06 2.585 2.055 2.585 2.055 2.605 1.82 2.605 1.82 2.465 2.055 2.465 2.055 2.525 2.06 2.525 ;
    END
  END SE
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0516 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.5925925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 23.287037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.165 0.92 1.09 0.92 1.09 1.14 1.12 1.14 1.12 1.2 1 1.2 1 1.14 1.03 1.14 1.03 0.72 1.165 0.72 ;
    END
  END SN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.695 2.61 3.215 2.61 3.215 2 3.345 2 3.345 1.89 3.595 1.89 3.595 2 3.695 2 ;
    END
  END ExtVDD
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.825 2.69 0.98 2.845 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.30535 LAYER Metal1 ;
    ANTENNADIFFAREA 3.9742 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2691 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.71516175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 145.1839465 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.56 2.83 5.525 2.83 5.525 3.135 5.465 3.135 5.465 2.83 5.43 2.83 5.43 2.495 5.465 2.495 5.465 2.07 5.525 2.07 5.525 2.495 5.56 2.495 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.30535 LAYER Metal1 ;
    ANTENNADIFFAREA 3.9742 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2691 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.71516175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 145.1839465 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.845 3.13 4.785 3.13 4.785 2.84 4.625 2.84 4.625 2.485 4.785 2.485 4.785 2.09 4.845 2.09 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 2.66 1.41 2.82 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.77 2.8 2.025 2.88 ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 3.48 0 3.48 0 3.36 0.85 3.36 0.85 2.97 0.91 2.97 0.91 3.36 1.3 3.36 1.3 2.94 1.36 2.94 1.36 3.36 1.92 3.36 1.92 2.94 1.98 2.94 1.98 3.36 3.215 3.36 3.215 3.025 3.275 3.025 3.275 3.36 3.635 3.36 3.635 3.025 3.695 3.025 3.695 3.36 4.99 3.36 4.99 2.87 5.05 2.87 5.05 3.36 5.67 3.36 5.67 2.875 5.73 2.875 5.73 3.36 6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6 0.06 5.265 0.06 5.265 0.35 5.26 0.35 5.26 0.465 5.2 0.465 5.2 0.32 5.205 0.32 5.205 0.06 3.79 0.06 3.79 0.465 3.73 0.465 3.73 0.06 0.95 0.06 0.95 0.32 1.185 0.32 1.185 0.44 1.125 0.44 1.125 0.465 0.89 0.465 0.89 0.06 0 0.06 0 -0.06 6 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.10185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.41 1.525 4.255 1.525 4.255 1.37 4.11 1.37 4.11 0.41 4.17 0.41 4.17 1.31 4.41 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.495 1.345 5.435 1.345 5.435 1.015 5.05 1.015 5.05 1.345 4.99 1.345 4.99 0.955 5.495 0.955 ;
      POLYGON 5.285 3.07 5.225 3.07 5.225 2.71 4.93 2.71 4.93 2.65 5.225 2.65 5.225 2.175 5.285 2.175 ;
      RECT 4.785 0.32 4.845 1.345 ;
      RECT 4.095 2.385 4.54 2.445 ;
      POLYGON 4.535 1.13 4.265 1.13 4.265 0.25 4.255 0.25 4.255 0.23 4.24 0.23 4.24 0.17 4.255 0.17 4.255 0.13 4.315 0.13 4.315 0.17 4.325 0.17 4.325 1.07 4.535 1.07 ;
      RECT 4.445 0.135 4.505 0.995 ;
      POLYGON 4.195 1.51 3.935 1.51 3.935 0.83 3.4 0.83 3.4 0.245 3.46 0.245 3.46 0.77 3.935 0.77 3.935 0.32 3.995 0.32 3.995 1.45 4.195 1.45 ;
      POLYGON 4.005 3.17 3.945 3.17 3.945 2.78 3.145 2.78 3.145 2.72 3.945 2.72 3.945 2 4.005 2 ;
      POLYGON 3.8 2.93 3.07 2.93 3.07 3.17 3.01 3.17 3.01 2 3.07 2 3.07 2.87 3.8 2.87 ;
      RECT 3.51 1.24 3.79 1.525 ;
      RECT 3.215 0.32 3.275 1.455 ;
      POLYGON 3.07 1.52 2.735 1.52 2.735 1.46 3.01 1.46 3.01 0.32 3.07 0.32 ;
      RECT 2.475 0.6 2.535 1.29 ;
      POLYGON 2.245 0.83 2.185 0.83 2.185 1.485 2.125 1.485 2.125 0.32 2.185 0.32 2.185 0.77 2.245 0.77 ;
      POLYGON 2.185 3.085 2.125 3.085 2.125 2.74 1.655 2.74 1.655 2.68 2.125 2.68 2.125 2.185 2.185 2.185 ;
      POLYGON 1.98 1.485 1.92 1.485 1.92 0.585 1.31 0.585 1.31 1.27 1.43 1.27 1.43 1.485 1.095 1.485 1.095 1.27 1.25 1.27 1.25 0.585 0.915 0.585 0.915 0.595 0.885 0.595 0.885 1.14 0.915 1.14 0.915 1.2 0.795 1.2 0.795 1.14 0.825 1.14 0.825 0.595 0.795 0.595 0.795 0.535 0.825 0.535 0.825 0.525 1.475 0.525 1.475 0.32 1.535 0.32 1.535 0.525 1.92 0.525 1.92 0.32 1.98 0.32 ;
      POLYGON 1.715 0.705 1.685 0.705 1.685 1.185 1.525 1.185 1.525 1.2 1.405 1.2 1.405 1.14 1.435 1.14 1.435 1.125 1.625 1.125 1.625 0.705 1.595 0.705 1.595 0.645 1.715 0.645 ;
      POLYGON 1.67 2.535 1.545 2.535 1.545 2.875 1.67 2.875 1.67 3.085 1.61 3.085 1.61 2.935 1.485 2.935 1.485 2.475 1.61 2.475 1.61 2.24 1.19 2.24 1.19 2.2 1.055 2.2 1.055 1.985 0.465 1.985 0.465 3.115 0.405 3.115 0.405 1.925 1.115 1.925 1.115 2.14 1.25 2.14 1.25 2.18 1.67 2.18 ;
      POLYGON 1.115 3.115 1.055 3.115 1.055 2.605 0.745 2.605 0.745 2.545 1.055 2.545 1.055 2.28 1.115 2.28 ;
      POLYGON 0.705 2.485 0.595 2.485 0.595 2.97 0.705 2.97 0.705 3.115 0.645 3.115 0.645 3.03 0.535 3.03 0.535 2.425 0.645 2.425 0.645 2.105 0.57 2.105 0.57 2.045 0.705 2.045 ;
      POLYGON 0.64 1.485 0.23 1.485 0.23 1.56 0.17 1.56 0.17 1.425 0.58 1.425 0.58 0.32 0.64 0.32 ;
      RECT 0.41 0.135 0.47 1.305 ;
      POLYGON 0.26 3.115 0.2 3.115 0.2 1.965 0.14 1.965 0.14 1.905 0.26 1.905 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END SRDFFNSX1

MACRO SRDFFNX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SRDFFNX1 0 0 ;
  SIZE 6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 1.77 5.73 1.77 5.73 2.46 5.67 2.46 5.67 1.77 5.05 1.77 5.05 2.48 4.99 2.48 4.99 1.77 1.98 1.77 1.98 2.4 1.92 2.4 1.92 1.77 1.33 1.77 1.33 2.08 1.27 2.08 1.27 1.77 -0.005 1.77 -0.005 1.65 0.89 1.65 0.89 1.27 0.95 1.27 0.95 1.65 5.23 1.65 5.23 1.13 5.29 1.13 5.29 1.65 6 1.65 ;
    END
  END VDD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.06 2.585 2.055 2.585 2.055 2.605 1.82 2.605 1.82 2.465 2.055 2.465 2.055 2.525 2.06 2.525 ;
    END
  END SE
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.695 2.61 3.215 2.61 3.215 2 3.345 2 3.345 1.89 3.595 1.89 3.595 2 3.695 2 ;
    END
  END ExtVDD
  PIN CKN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.8 2.69 0.985 2.825 ;
    END
  END CKN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1058 LAYER Metal1 ;
    ANTENNADIFFAREA 3.822325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2691 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.97361575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 139.8996655 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.565 2.825 5.525 2.825 5.525 3.135 5.465 3.135 5.465 2.825 5.435 2.825 5.435 2.495 5.465 2.495 5.465 2.07 5.525 2.07 5.525 2.495 5.565 2.495 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1058 LAYER Metal1 ;
    ANTENNADIFFAREA 3.822325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2691 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.97361575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 139.8996655 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.845 3.13 4.785 3.13 4.785 2.84 4.625 2.84 4.625 2.48 4.785 2.48 4.785 2.09 4.845 2.09 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.235 2.66 1.41 2.82 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.111111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.775 2.8 2.025 2.88 ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 3.48 0 3.48 0 3.36 0.85 3.36 0.85 2.97 0.91 2.97 0.91 3.36 1.3 3.36 1.3 2.94 1.36 2.94 1.36 3.36 1.92 3.36 1.92 2.94 1.98 2.94 1.98 3.36 3.215 3.36 3.215 3.025 3.275 3.025 3.275 3.36 3.635 3.36 3.635 3.025 3.695 3.025 3.695 3.36 4.99 3.36 4.99 2.87 5.05 2.87 5.05 3.36 5.67 3.36 5.67 2.875 5.73 2.875 5.73 3.36 6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6 0.06 5.155 0.06 5.155 0.465 5.095 0.465 5.095 0.06 3.79 0.06 3.79 0.465 3.73 0.465 3.73 0.06 0.95 0.06 0.95 0.465 0.89 0.465 0.89 0.06 0 0.06 0 -0.06 6 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.10185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.41 1.525 4.255 1.525 4.255 1.37 4.11 1.37 4.11 0.41 4.17 0.41 4.17 1.31 4.41 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.495 1.345 5.435 1.345 5.435 1.015 5.05 1.015 5.05 1.345 4.99 1.345 4.99 0.955 5.495 0.955 ;
      POLYGON 5.285 3.07 5.225 3.07 5.225 2.71 4.93 2.71 4.93 2.65 5.225 2.65 5.225 2.175 5.285 2.175 ;
      RECT 4.785 0.32 4.845 1.345 ;
      RECT 4.095 2.385 4.54 2.445 ;
      POLYGON 4.535 1.07 4.265 1.07 4.265 0.25 4.255 0.25 4.255 0.23 4.24 0.23 4.24 0.17 4.255 0.17 4.255 0.13 4.315 0.13 4.315 0.17 4.325 0.17 4.325 1.01 4.535 1.01 ;
      POLYGON 4.195 1.51 3.935 1.51 3.935 0.83 3.4 0.83 3.4 0.245 3.46 0.245 3.46 0.77 3.935 0.77 3.935 0.32 3.995 0.32 3.995 1.45 4.195 1.45 ;
      POLYGON 4.005 3.17 3.945 3.17 3.945 2.78 3.145 2.78 3.145 2.72 3.945 2.72 3.945 2 4.005 2 ;
      POLYGON 3.8 2.93 3.07 2.93 3.07 3.17 3.01 3.17 3.01 2 3.07 2 3.07 2.87 3.8 2.87 ;
      RECT 3.51 1.24 3.79 1.525 ;
      RECT 3.215 0.32 3.275 1.455 ;
      POLYGON 3.07 1.52 2.735 1.52 2.735 1.46 3.01 1.46 3.01 0.32 3.07 0.32 ;
      RECT 2.475 0.6 2.535 1.29 ;
      POLYGON 2.245 0.83 2.185 0.83 2.185 1.485 2.125 1.485 2.125 0.32 2.185 0.32 2.185 0.77 2.245 0.77 ;
      POLYGON 2.185 3.085 2.125 3.085 2.125 2.74 1.655 2.74 1.655 2.68 2.125 2.68 2.125 2.185 2.185 2.185 ;
      POLYGON 1.98 1.485 1.92 1.485 1.92 0.585 1.155 0.585 1.155 1.485 1.095 1.485 1.095 0.585 0.915 0.585 0.915 0.595 0.885 0.595 0.885 1.14 0.915 1.14 0.915 1.2 0.795 1.2 0.795 1.14 0.825 1.14 0.825 0.595 0.795 0.595 0.795 0.535 0.825 0.535 0.825 0.525 1.095 0.525 1.095 0.32 1.155 0.32 1.155 0.525 1.92 0.525 1.92 0.32 1.98 0.32 ;
      POLYGON 1.67 2.535 1.545 2.535 1.545 2.875 1.67 2.875 1.67 3.085 1.61 3.085 1.61 2.935 1.485 2.935 1.485 2.475 1.61 2.475 1.61 2.24 1.19 2.24 1.19 2.2 1.055 2.2 1.055 1.985 0.465 1.985 0.465 3.115 0.405 3.115 0.405 1.925 1.115 1.925 1.115 2.14 1.25 2.14 1.25 2.18 1.67 2.18 ;
      POLYGON 1.115 3.115 1.055 3.115 1.055 2.605 0.745 2.605 0.745 2.545 1.055 2.545 1.055 2.28 1.115 2.28 ;
      POLYGON 0.705 2.49 0.595 2.49 0.595 2.97 0.705 2.97 0.705 3.115 0.645 3.115 0.645 3.03 0.535 3.03 0.535 2.43 0.645 2.43 0.645 2.105 0.57 2.105 0.57 2.045 0.705 2.045 ;
      POLYGON 0.64 1.485 0.23 1.485 0.23 1.56 0.17 1.56 0.17 1.425 0.58 1.425 0.58 0.32 0.64 0.32 ;
      RECT 0.41 0.135 0.47 1.305 ;
      POLYGON 0.26 3.115 0.2 3.115 0.2 1.965 0.14 1.965 0.14 1.905 0.26 1.905 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END SRDFFNX1

MACRO SRDFFQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SRDFFQX1 0 0 ;
  SIZE 5.8 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.8 1.77 5.31 1.77 5.31 2.46 5.25 2.46 5.25 1.77 1.985 1.77 1.985 2.4 1.925 2.4 1.925 1.77 1.335 1.77 1.335 2.08 1.275 2.08 1.275 1.77 0 1.77 0 1.65 0.895 1.65 0.895 1.27 0.955 1.27 0.955 1.65 1.05 1.65 1.05 1.485 1.11 1.485 1.11 1.65 1.46 1.65 1.46 1.27 1.52 1.27 1.52 1.65 5.34 1.65 5.34 1.13 5.4 1.13 5.4 1.65 5.8 1.65 ;
    END
  END VDD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.065 2.585 2.06 2.585 2.06 2.605 1.825 2.605 1.825 2.465 2.06 2.465 2.06 2.525 2.065 2.525 ;
    END
  END SE
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        RECT 3.22 2 3.7 2.61 ;
    END
  END ExtVDD
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.961525 LAYER Metal1 ;
    ANTENNADIFFAREA 3.423225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.22365 LAYER Metal1 ;
      ANTENNAMAXAREACAR 22.18432825 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 168.169014 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 5.045 2.07 5.105 3.135 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.22 2.66 1.415 2.79 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.755 2.8 2.05 2.87 ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.86 3.48 0 3.48 0 3.36 0.855 3.36 0.855 2.97 0.915 2.97 0.915 3.36 1.305 3.36 1.305 2.94 1.365 2.94 1.365 3.36 1.925 3.36 1.925 2.96 1.985 2.96 1.985 3.36 3.22 3.36 3.22 3.025 3.28 3.025 3.28 3.36 3.64 3.36 3.64 3.025 3.7 3.025 3.7 3.36 5.25 3.36 5.25 2.875 5.31 2.875 5.31 3.36 5.86 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.86 0.06 5.605 0.06 5.605 0.465 5.545 0.465 5.545 0.06 3.755 0.06 3.755 0.34 3.695 0.34 3.695 0.06 1.315 0.06 1.315 0.465 1.255 0.465 1.255 0.06 0.955 0.06 0.955 0.465 0.895 0.465 0.895 0.06 0 0.06 0 -0.06 5.86 -0.06 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.85185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.725 2.565 0.985 2.675 ;
    END
  END CK
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.26 1.095 4.5 1.235 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.605 1.345 5.545 1.345 5.545 1.015 5.055 1.015 5.055 1.345 4.995 1.345 4.995 0.955 5.605 0.955 ;
      POLYGON 5.4 0.545 4.995 0.545 4.995 0.32 5.055 0.32 5.055 0.485 5.34 0.485 5.34 0.32 5.4 0.32 ;
      POLYGON 4.85 1.345 4.79 1.345 4.79 0.425 4.575 0.425 4.575 0.365 4.79 0.365 4.79 0.32 4.85 0.32 ;
      POLYGON 4.705 0.665 4.645 0.665 4.645 1.375 2.58 1.375 2.58 1.315 4.585 1.315 4.585 0.51 4.675 0.51 4.675 0.605 4.705 0.605 ;
      RECT 4.1 2.615 4.545 2.675 ;
      POLYGON 4.515 1 4.27 1 4.27 0.25 4.26 0.25 4.26 0.23 4.245 0.23 4.245 0.17 4.26 0.17 4.26 0.13 4.32 0.13 4.32 0.17 4.33 0.17 4.33 0.94 4.515 0.94 ;
      POLYGON 4.2 1.22 4 1.22 4 1.255 3.94 1.255 3.94 1.13 4 1.13 4 1.16 4.14 1.16 4.14 0.415 4 0.415 4 0.47 3.515 0.47 3.515 0.3 3.4 0.3 3.4 0.24 3.575 0.24 3.575 0.41 3.94 0.41 3.94 0.32 4 0.32 4 0.355 4.2 0.355 ;
      POLYGON 4.07 0.615 3.535 0.615 3.535 0.65 3.415 0.65 3.415 0.59 3.475 0.59 3.475 0.555 4.07 0.555 ;
      POLYGON 4.01 3.17 3.95 3.17 3.95 2.78 3.15 2.78 3.15 2.72 3.95 2.72 3.95 2 4.01 2 ;
      POLYGON 3.805 2.93 3.075 2.93 3.075 3.17 3.015 3.17 3.015 2 3.075 2 3.075 2.87 3.805 2.87 ;
      RECT 3.54 1.13 3.795 1.25 ;
      POLYGON 3.455 1.25 3.22 1.25 3.22 0.32 3.28 0.32 3.28 1.19 3.395 1.19 3.395 1.13 3.455 1.13 ;
      POLYGON 3.075 1.255 3.015 1.255 3.015 0.65 2.19 0.65 2.19 1.485 2.13 1.485 2.13 0.32 2.19 0.32 2.19 0.59 2.955 0.59 2.955 0.58 3.015 0.58 3.015 0.32 3.075 0.32 ;
      POLYGON 2.235 3.035 2.1 3.035 2.1 2.975 2.175 2.975 2.175 2.74 1.66 2.74 1.66 2.68 2.175 2.68 2.175 2.4 2.13 2.4 2.13 2.185 2.235 2.185 ;
      POLYGON 1.985 1.485 1.925 1.485 1.925 0.585 1.315 0.585 1.315 1.485 1.255 1.485 1.255 0.585 0.92 0.585 0.92 0.595 0.89 0.595 0.89 1.14 0.92 1.14 0.92 1.2 0.8 1.2 0.8 1.14 0.83 1.14 0.83 0.595 0.8 0.595 0.8 0.535 0.83 0.535 0.83 0.525 1.46 0.525 1.46 0.32 1.52 0.32 1.52 0.525 1.925 0.525 1.925 0.32 1.985 0.32 ;
      POLYGON 1.675 2.535 1.55 2.535 1.55 2.875 1.675 2.875 1.675 3.085 1.615 3.085 1.615 2.935 1.49 2.935 1.49 2.475 1.615 2.475 1.615 2.24 1.195 2.24 1.195 2.2 1.06 2.2 1.06 1.985 0.47 1.985 0.47 3.115 0.41 3.115 0.41 1.925 1.12 1.925 1.12 2.14 1.255 2.14 1.255 2.18 1.675 2.18 ;
      POLYGON 1.12 3.115 1.06 3.115 1.06 2.795 0.75 2.795 0.75 2.735 1.06 2.735 1.06 2.28 1.12 2.28 ;
      POLYGON 0.71 2.5 0.645 2.5 0.645 2.97 0.71 2.97 0.71 3.115 0.65 3.115 0.65 3.03 0.585 3.03 0.585 2.44 0.65 2.44 0.65 2.18 0.71 2.18 ;
      POLYGON 0.645 1.485 0.235 1.485 0.235 1.56 0.175 1.56 0.175 1.425 0.585 1.425 0.585 0.32 0.645 0.32 ;
      RECT 0.415 0.135 0.475 1.305 ;
      POLYGON 0.265 3.115 0.205 3.115 0.205 1.965 0.145 1.965 0.145 1.905 0.265 1.905 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END SRDFFQX1

MACRO SRDFFRQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SRDFFRQX1 0 0 ;
  SIZE 5.6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 5.445 1.77 5.445 2.46 5.385 2.46 5.385 1.77 2.18 1.77 2.18 2.4 2.12 2.4 2.12 1.77 1.53 1.77 1.53 2.08 1.47 2.08 1.47 1.77 0 1.77 0 1.65 0.245 1.65 0.245 1.05 0.305 1.05 0.305 1.65 1.09 1.65 1.09 1.27 1.15 1.27 1.15 1.65 1.64 1.65 1.64 1.27 1.7 1.27 1.7 1.65 5.4 1.65 5.4 1.13 5.46 1.13 5.46 1.65 5.6 1.65 ;
    END
  END VDD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.26 2.585 2.255 2.585 2.255 2.605 2.02 2.605 2.02 2.465 2.255 2.465 2.255 2.525 2.26 2.525 ;
    END
  END SE
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.895 2.61 3.415 2.61 3.415 2 3.545 2 3.545 1.89 3.795 1.89 3.795 2 3.895 2 ;
    END
  END ExtVDD
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.385 0.905 0.375 0.905 0.375 0.98 0.245 0.98 0.245 0.74 0.375 0.74 0.375 0.845 0.385 0.845 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.937475 LAYER Metal1 ;
    ANTENNADIFFAREA 3.641925 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.25605 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.2832455 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 145.14352675 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.24 3.135 5.18 3.135 5.18 2.845 5.015 2.845 5.015 2.685 5.18 2.685 5.18 2.07 5.24 2.07 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.9444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.415 2.66 1.61 2.84 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.97 2.8 2.225 2.88 ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 3.48 0 3.48 0 3.36 1.05 3.36 1.05 2.97 1.11 2.97 1.11 3.36 1.5 3.36 1.5 2.94 1.56 2.94 1.56 3.36 2.12 3.36 2.12 2.94 2.18 2.94 2.18 3.36 3.415 3.36 3.415 3.025 3.475 3.025 3.475 3.36 3.835 3.36 3.835 3.025 3.895 3.025 3.895 3.36 5.385 3.36 5.385 2.875 5.445 2.875 5.445 3.36 5.6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5.255 0.06 5.255 0.32 5.26 0.32 5.26 0.465 5.2 0.465 5.2 0.35 5.195 0.35 5.195 0.06 3.99 0.06 3.99 0.465 3.93 0.465 3.93 0.06 1.56 0.06 1.56 0.465 1.5 0.465 1.5 0.06 1.15 0.06 1.15 0.465 1.09 0.465 1.09 0.06 0.305 0.06 0.305 0.465 0.245 0.465 0.245 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
  END VSS
  PIN CK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.025 2.69 1.18 2.845 ;
    END
  END CK
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.10185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.61 1.525 4.455 1.525 4.455 1.37 4.31 1.37 4.31 0.41 4.37 0.41 4.37 1.31 4.61 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.465 0.625 4.99 0.625 4.99 0.32 5.055 0.32 5.055 0.465 5.05 0.465 5.05 0.565 5.405 0.565 5.405 0.29 5.465 0.29 ;
      POLYGON 5.045 1.345 4.985 1.345 4.985 0.83 4.85 0.83 4.85 0.86 4.79 0.86 4.79 0.32 4.85 0.32 4.85 0.77 5.045 0.77 ;
      RECT 4.295 2.385 4.785 2.445 ;
      POLYGON 4.78 1.235 4.465 1.235 4.465 0.25 4.455 0.25 4.455 0.23 4.44 0.23 4.44 0.17 4.455 0.17 4.455 0.13 4.515 0.13 4.515 0.17 4.525 0.17 4.525 1.175 4.78 1.175 ;
      RECT 4.66 0.13 4.72 1.075 ;
      POLYGON 4.395 1.51 4.135 1.51 4.135 0.83 3.6 0.83 3.6 0.245 3.66 0.245 3.66 0.77 4.135 0.77 4.135 0.32 4.195 0.32 4.195 1.45 4.395 1.45 ;
      POLYGON 4.205 3.17 4.145 3.17 4.145 2.78 3.345 2.78 3.345 2.72 4.145 2.72 4.145 2 4.205 2 ;
      POLYGON 4 2.93 3.27 2.93 3.27 3.17 3.21 3.17 3.21 2 3.27 2 3.27 2.87 4 2.87 ;
      RECT 3.71 1.24 3.99 1.525 ;
      RECT 3.415 0.32 3.475 1.455 ;
      POLYGON 3.27 1.52 2.935 1.52 2.935 1.46 3.21 1.46 3.21 0.32 3.27 0.32 ;
      RECT 2.675 0.6 2.735 1.29 ;
      POLYGON 2.445 0.83 2.385 0.83 2.385 1.485 2.325 1.485 2.325 0.32 2.385 0.32 2.385 0.77 2.445 0.77 ;
      POLYGON 2.385 3.085 2.325 3.085 2.325 2.74 1.855 2.74 1.855 2.68 2.325 2.68 2.325 2.185 2.385 2.185 ;
      POLYGON 2.18 1.485 2.12 1.485 2.12 0.585 1.39 0.585 1.39 1.485 1.33 1.485 1.33 0.585 1.115 0.585 1.115 0.595 1.085 0.595 1.085 1.14 1.115 1.14 1.115 1.2 0.995 1.2 0.995 1.14 1.025 1.14 1.025 0.595 0.995 0.595 0.995 0.535 1.025 0.535 1.025 0.525 1.295 0.525 1.295 0.32 1.355 0.32 1.355 0.525 2.12 0.525 2.12 0.32 2.18 0.32 ;
      POLYGON 1.87 2.535 1.745 2.535 1.745 2.875 1.87 2.875 1.87 3.085 1.81 3.085 1.81 2.935 1.685 2.935 1.685 2.475 1.81 2.475 1.81 2.24 1.39 2.24 1.39 2.2 1.255 2.2 1.255 1.95 0.665 1.95 0.665 3.115 0.605 3.115 0.605 1.89 1.315 1.89 1.315 2.14 1.45 2.14 1.45 2.18 1.87 2.18 ;
      POLYGON 1.315 3.115 1.255 3.115 1.255 2.605 0.975 2.605 0.975 2.545 1.255 2.545 1.255 2.28 1.315 2.28 ;
      POLYGON 0.905 3.115 0.845 3.115 0.845 2.105 0.735 2.105 0.735 2.045 0.905 2.045 ;
      POLYGON 0.84 1.485 0.43 1.485 0.43 1.56 0.37 1.56 0.37 1.425 0.78 1.425 0.78 0.32 0.84 0.32 ;
      RECT 0.61 0.135 0.67 1.305 ;
      POLYGON 0.55 0.985 0.51 0.985 0.51 1.265 0.45 1.265 0.45 0.32 0.51 0.32 0.51 0.865 0.55 0.865 ;
      POLYGON 0.46 3.115 0.4 3.115 0.4 1.965 0.34 1.965 0.34 1.905 0.46 1.905 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END SRDFFRQX1

MACRO SRDFFRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SRDFFRX1 0 0 ;
  SIZE 6.2 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 5.93 1.77 5.93 2.46 5.87 2.46 5.87 1.77 5.25 1.77 5.25 2.48 5.19 2.48 5.19 1.77 2.18 1.77 2.18 2.4 2.12 2.4 2.12 1.77 1.53 1.77 1.53 2.08 1.47 2.08 1.47 1.77 -0.005 1.77 -0.005 1.65 0.245 1.65 0.245 1.05 0.305 1.05 0.305 1.65 1.09 1.65 1.09 1.27 1.15 1.27 1.15 1.65 1.745 1.65 1.745 1.27 1.805 1.27 1.805 1.65 5.43 1.65 5.43 1.13 5.49 1.13 5.49 1.65 6.2 1.65 ;
    END
  END VDD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.26 2.585 2.255 2.585 2.255 2.605 2.02 2.605 2.02 2.465 2.255 2.465 2.255 2.525 2.26 2.525 ;
    END
  END SE
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.895 2.61 3.415 2.61 3.415 2 3.545 2 3.545 1.89 3.795 1.89 3.795 2 3.895 2 ;
    END
  END ExtVDD
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.385 0.905 0.375 0.905 0.375 0.98 0.245 0.98 0.245 0.74 0.375 0.74 0.375 0.845 0.385 0.845 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.45605 LAYER Metal1 ;
    ANTENNADIFFAREA 4.111775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3015 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.0963515 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 135.43283575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.77 2.83 5.725 2.83 5.725 3.135 5.665 3.135 5.665 2.83 5.625 2.83 5.625 2.5 5.665 2.5 5.665 2.07 5.725 2.07 5.725 2.5 5.77 2.5 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.45605 LAYER Metal1 ;
    ANTENNADIFFAREA 4.111775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3015 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.0963515 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 135.43283575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.045 3.13 4.985 3.13 4.985 2.845 4.825 2.845 4.825 2.485 4.985 2.485 4.985 2.09 5.045 2.09 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.435 2.66 1.61 2.82 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.388889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.965 2.8 2.23 2.88 ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 3.48 0 3.48 0 3.36 1.05 3.36 1.05 2.97 1.11 2.97 1.11 3.36 1.5 3.36 1.5 2.94 1.56 2.94 1.56 3.36 2.12 3.36 2.12 2.94 2.18 2.94 2.18 3.36 3.415 3.36 3.415 3.025 3.475 3.025 3.475 3.36 3.835 3.36 3.835 3.025 3.895 3.025 3.895 3.36 5.19 3.36 5.19 2.87 5.25 2.87 5.25 3.36 5.87 3.36 5.87 2.875 5.93 2.875 5.93 3.36 6.2 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 5.86 0.06 5.86 0.465 5.8 0.465 5.8 0.06 5.45 0.06 5.45 0.465 5.39 0.465 5.39 0.06 3.99 0.06 3.99 0.465 3.93 0.465 3.93 0.06 1.84 0.06 1.84 0.465 1.78 0.465 1.78 0.06 1.15 0.06 1.15 0.465 1.09 0.465 1.09 0.06 0.305 0.06 0.305 0.465 0.245 0.465 0.245 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.025 2.69 1.18 2.845 ;
    END
  END CK
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.10185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.61 1.525 4.455 1.525 4.455 1.37 4.31 1.37 4.31 0.41 4.37 0.41 4.37 1.31 4.61 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.8 1.345 5.74 1.345 5.74 1.015 5.25 1.015 5.25 1.345 5.19 1.345 5.19 0.955 5.8 0.955 ;
      POLYGON 5.655 0.67 5.19 0.67 5.19 0.32 5.25 0.32 5.25 0.61 5.595 0.61 5.595 0.32 5.655 0.32 ;
      POLYGON 5.485 3.07 5.425 3.07 5.425 2.71 5.13 2.71 5.13 2.65 5.425 2.65 5.425 2.175 5.485 2.175 ;
      RECT 4.985 0.32 5.045 1.345 ;
      POLYGON 4.81 1.07 4.465 1.07 4.465 0.25 4.455 0.25 4.455 0.23 4.44 0.23 4.44 0.17 4.455 0.17 4.455 0.13 4.515 0.13 4.515 0.17 4.525 0.17 4.525 1.01 4.81 1.01 ;
      RECT 4.295 2.385 4.74 2.445 ;
      POLYGON 4.395 1.51 4.135 1.51 4.135 0.83 3.6 0.83 3.6 0.245 3.66 0.245 3.66 0.77 4.135 0.77 4.135 0.32 4.195 0.32 4.195 1.45 4.395 1.45 ;
      POLYGON 4.205 3.17 4.145 3.17 4.145 2.78 3.345 2.78 3.345 2.72 4.145 2.72 4.145 2 4.205 2 ;
      POLYGON 4 2.93 3.27 2.93 3.27 3.17 3.21 3.17 3.21 2 3.27 2 3.27 2.87 4 2.87 ;
      RECT 3.71 1.24 3.99 1.525 ;
      RECT 3.415 0.32 3.475 1.455 ;
      POLYGON 3.27 1.52 2.935 1.52 2.935 1.46 3.21 1.46 3.21 0.32 3.27 0.32 ;
      RECT 2.675 0.6 2.735 1.29 ;
      POLYGON 2.385 3.085 2.325 3.085 2.325 2.74 1.855 2.74 1.855 2.68 2.325 2.68 2.325 2.185 2.385 2.185 ;
      POLYGON 2.31 0.83 2.25 0.83 2.25 1.485 2.19 1.485 2.19 0.32 2.25 0.32 2.25 0.77 2.31 0.77 ;
      POLYGON 2.045 1.485 1.985 1.485 1.985 0.585 1.495 0.585 1.495 1.485 1.435 1.485 1.435 0.585 1.115 0.585 1.115 0.595 1.085 0.595 1.085 1.14 1.115 1.14 1.115 1.2 0.995 1.2 0.995 1.14 1.025 1.14 1.025 0.595 0.995 0.595 0.995 0.535 1.025 0.535 1.025 0.525 1.295 0.525 1.295 0.32 1.355 0.32 1.355 0.525 1.985 0.525 1.985 0.32 2.045 0.32 ;
      POLYGON 1.87 2.535 1.745 2.535 1.745 2.875 1.87 2.875 1.87 3.085 1.81 3.085 1.81 2.935 1.685 2.935 1.685 2.475 1.81 2.475 1.81 2.24 1.39 2.24 1.39 2.2 1.255 2.2 1.255 1.955 0.665 1.955 0.665 3.115 0.605 3.115 0.605 1.895 1.315 1.895 1.315 2.14 1.45 2.14 1.45 2.18 1.87 2.18 ;
      POLYGON 1.315 3.115 1.255 3.115 1.255 2.605 0.97 2.605 0.97 2.545 1.255 2.545 1.255 2.28 1.315 2.28 ;
      RECT 1.19 0.68 1.25 1.09 ;
      POLYGON 0.905 3.115 0.845 3.115 0.845 2.115 0.74 2.115 0.74 2.055 0.905 2.055 ;
      POLYGON 0.84 1.485 0.43 1.485 0.43 1.56 0.37 1.56 0.37 1.425 0.78 1.425 0.78 0.32 0.84 0.32 ;
      RECT 0.61 0.135 0.67 1.305 ;
      POLYGON 0.55 0.95 0.51 0.95 0.51 1.265 0.45 1.265 0.45 0.32 0.51 0.32 0.51 0.83 0.55 0.83 ;
      POLYGON 0.46 3.115 0.4 3.115 0.4 1.965 0.34 1.965 0.34 1.905 0.46 1.905 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END SRDFFRX1

MACRO SRDFFSQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SRDFFSQX1 0 0 ;
  SIZE 6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 1.77 5.625 1.77 5.625 2.46 5.565 2.46 5.565 1.77 1.98 1.77 1.98 2.4 1.92 2.4 1.92 1.77 1.33 1.77 1.33 2.08 1.27 2.08 1.27 1.77 -0.005 1.77 -0.005 1.65 0.89 1.65 0.89 1.27 0.95 1.27 0.95 1.65 1.045 1.65 1.045 1.27 1.105 1.27 1.105 1.65 1.455 1.65 1.455 1.27 1.515 1.27 1.515 1.65 5.23 1.65 5.23 1.13 5.29 1.13 5.29 1.65 5.64 1.65 5.64 1.13 5.7 1.13 5.7 1.65 6 1.65 ;
    END
  END VDD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.06 2.585 2.055 2.585 2.055 2.605 1.82 2.605 1.82 2.465 2.055 2.465 2.055 2.525 2.06 2.525 ;
    END
  END SE
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0516 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.5925925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 23.37962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.17 0.94 1.105 0.94 1.105 1.14 1.135 1.14 1.135 1.2 1.015 1.2 1.015 1.14 1.045 1.14 1.045 0.94 1.025 0.94 1.025 0.72 1.17 0.72 ;
    END
  END SN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.695 2.61 3.215 2.61 3.215 2 3.345 2 3.345 1.89 3.595 1.89 3.595 2 3.695 2 ;
    END
  END ExtVDD
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.991975 LAYER Metal1 ;
    ANTENNADIFFAREA 3.716825 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.22365 LAYER Metal1 ;
      ANTENNAMAXAREACAR 22.3204785 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 163.715627 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.42 3.135 5.36 3.135 5.36 2.835 5.225 2.835 5.225 2.495 5.36 2.495 5.36 2.07 5.42 2.07 ;
    END
  END Q
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.12962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.775 2.665 0.98 2.845 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 2.66 1.41 2.79 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.75 2.8 2.045 2.87 ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 3.48 0 3.48 0 3.36 0.85 3.36 0.85 2.97 0.91 2.97 0.91 3.36 1.3 3.36 1.3 2.94 1.36 2.94 1.36 3.36 1.92 3.36 1.92 2.94 1.98 2.94 1.98 3.36 3.215 3.36 3.215 3.025 3.275 3.025 3.275 3.36 3.635 3.36 3.635 3.025 3.695 3.025 3.695 3.36 5.565 3.36 5.565 2.875 5.625 2.875 5.625 3.36 6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6 0.06 5.265 0.06 5.265 0.35 5.26 0.35 5.26 0.465 5.2 0.465 5.2 0.32 5.205 0.32 5.205 0.06 3.79 0.06 3.79 0.465 3.73 0.465 3.73 0.06 0.95 0.06 0.95 0.32 1.125 0.32 1.125 0.465 0.89 0.465 0.89 0.06 0 0.06 0 -0.06 6 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.10185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.41 1.525 4.255 1.525 4.255 1.37 4.11 1.37 4.11 0.41 4.17 0.41 4.17 1.31 4.41 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.495 1.345 5.435 1.345 5.435 1.015 5.05 1.015 5.05 1.345 4.99 1.345 4.99 0.955 5.495 0.955 ;
      RECT 4.785 0.32 4.845 1.345 ;
      RECT 4.095 2.385 4.54 2.445 ;
      POLYGON 4.535 1.13 4.265 1.13 4.265 0.25 4.255 0.25 4.255 0.23 4.24 0.23 4.24 0.17 4.255 0.17 4.255 0.13 4.315 0.13 4.315 0.17 4.325 0.17 4.325 1.07 4.535 1.07 ;
      RECT 4.445 0.135 4.505 0.995 ;
      POLYGON 4.195 1.51 3.935 1.51 3.935 0.83 3.4 0.83 3.4 0.245 3.46 0.245 3.46 0.77 3.935 0.77 3.935 0.32 3.995 0.32 3.995 1.45 4.195 1.45 ;
      POLYGON 4.005 3.17 3.945 3.17 3.945 2.78 3.145 2.78 3.145 2.72 3.945 2.72 3.945 2 4.005 2 ;
      POLYGON 3.8 2.93 3.07 2.93 3.07 3.17 3.01 3.17 3.01 2 3.07 2 3.07 2.87 3.8 2.87 ;
      RECT 3.51 1.24 3.79 1.525 ;
      RECT 3.215 0.32 3.275 1.455 ;
      POLYGON 3.07 1.52 2.735 1.52 2.735 1.46 3.01 1.46 3.01 0.32 3.07 0.32 ;
      RECT 2.475 0.6 2.535 1.29 ;
      POLYGON 2.245 0.83 2.185 0.83 2.185 1.485 2.125 1.485 2.125 0.32 2.185 0.32 2.185 0.77 2.245 0.77 ;
      POLYGON 2.185 3.085 2.125 3.085 2.125 2.74 1.655 2.74 1.655 2.68 2.125 2.68 2.125 2.185 2.185 2.185 ;
      POLYGON 1.98 1.485 1.92 1.485 1.92 0.585 1.31 0.585 1.31 1.485 1.25 1.485 1.25 0.585 0.915 0.585 0.915 0.595 0.885 0.595 0.885 1.14 0.915 1.14 0.915 1.2 0.795 1.2 0.795 1.14 0.825 1.14 0.825 0.595 0.795 0.595 0.795 0.535 0.825 0.535 0.825 0.525 1.375 0.525 1.375 0.32 1.435 0.32 1.435 0.525 1.92 0.525 1.92 0.32 1.98 0.32 ;
      POLYGON 1.67 2.535 1.545 2.535 1.545 2.875 1.67 2.875 1.67 3.085 1.61 3.085 1.61 2.935 1.485 2.935 1.485 2.475 1.61 2.475 1.61 2.21 1.145 2.21 1.145 2.18 1.055 2.18 1.055 1.93 0.465 1.93 0.465 3.115 0.405 3.115 0.405 1.87 1.115 1.87 1.115 2.12 1.205 2.12 1.205 2.15 1.67 2.15 ;
      RECT 1.38 0.67 1.44 1.13 ;
      POLYGON 1.115 3.115 1.055 3.115 1.055 2.56 0.775 2.56 0.775 2.5 1.055 2.5 1.055 2.28 1.115 2.28 ;
      POLYGON 0.705 3.115 0.645 3.115 0.645 2.105 0.58 2.105 0.58 2.1 0.55 2.1 0.55 2.04 0.67 2.04 0.67 2.045 0.705 2.045 ;
      POLYGON 0.64 1.485 0.23 1.485 0.23 1.56 0.17 1.56 0.17 1.425 0.58 1.425 0.58 0.32 0.64 0.32 ;
      RECT 0.41 0.135 0.47 1.305 ;
      POLYGON 0.26 3.115 0.2 3.115 0.2 1.965 0.14 1.965 0.14 1.905 0.26 1.905 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END SRDFFSQX1

MACRO SRDFFSRQX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SRDFFSRQX1 0 0 ;
  SIZE 6.2 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 5.93 1.77 5.93 2.46 5.87 2.46 5.87 1.77 2.18 1.77 2.18 2.4 2.12 2.4 2.12 1.77 1.53 1.77 1.53 2.08 1.47 2.08 1.47 1.77 -0.005 1.77 -0.005 1.65 0.245 1.65 0.245 1.05 0.305 1.05 0.305 1.65 1.09 1.65 1.09 1.27 1.15 1.27 1.15 1.65 1.88 1.65 1.88 1.27 1.94 1.27 1.94 1.65 5.43 1.65 5.43 1.13 5.49 1.13 5.49 1.65 5.945 1.65 5.945 1.13 6.005 1.13 6.005 1.65 6.2 1.65 ;
    END
  END VDD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.26 2.585 2.255 2.585 2.255 2.605 2.02 2.605 2.02 2.465 2.255 2.465 2.255 2.525 2.26 2.525 ;
    END
  END SE
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0516 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.5925925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 23.47222225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 0.92 1.29 0.92 1.29 1.14 1.32 1.14 1.32 1.2 1.2 1.2 1.2 1.14 1.23 1.14 1.23 0.92 1.21 0.92 1.21 0.72 1.365 0.72 ;
    END
  END SN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.895 2.61 3.415 2.61 3.415 2 3.545 2 3.545 1.89 3.795 1.89 3.795 2 3.895 2 ;
    END
  END ExtVDD
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.9444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.385 0.905 0.375 0.905 0.375 0.98 0.25 0.98 0.25 0.74 0.375 0.74 0.375 0.845 0.385 0.845 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.4432 LAYER Metal1 ;
    ANTENNADIFFAREA 3.9912 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.25605 LAYER Metal1 ;
      ANTENNAMAXAREACAR 21.258348 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 158.8166375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.765 2.825 5.725 2.825 5.725 3.135 5.665 3.135 5.665 2.825 5.63 2.825 5.63 2.5 5.665 2.5 5.665 2.07 5.725 2.07 5.725 2.5 5.765 2.5 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.415 2.66 1.61 2.82 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.95 2.8 2.245 2.87 ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 3.48 0 3.48 0 3.36 1.05 3.36 1.05 2.97 1.11 2.97 1.11 3.36 1.5 3.36 1.5 2.94 1.56 2.94 1.56 3.36 2.12 3.36 2.12 2.94 2.18 2.94 2.18 3.36 3.415 3.36 3.415 3.025 3.475 3.025 3.475 3.36 3.835 3.36 3.835 3.025 3.895 3.025 3.895 3.36 5.87 3.36 5.87 2.875 5.93 2.875 5.93 3.36 6.2 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 6.065 0.06 6.065 0.465 6.005 0.465 6.005 0.06 3.99 0.06 3.99 0.465 3.93 0.465 3.93 0.06 1.15 0.06 1.15 0.32 1.325 0.32 1.325 0.465 1.09 0.465 1.09 0.06 0.305 0.06 0.305 0.465 0.245 0.465 0.245 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.10185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.61 1.525 4.455 1.525 4.455 1.37 4.31 1.37 4.31 0.41 4.37 0.41 4.37 1.31 4.61 1.31 ;
    END
  END RT
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.85185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.975 2.69 1.18 2.855 ;
    END
  END CK
  OBS
    LAYER Metal1 ;
      POLYGON 5.86 0.465 5.8 0.465 5.8 0.26 5.45 0.26 5.45 0.465 5.39 0.465 5.39 0.2 5.86 0.2 ;
      POLYGON 5.8 1.345 5.74 1.345 5.74 1.015 5.25 1.015 5.25 1.345 5.19 1.345 5.19 0.955 5.8 0.955 ;
      POLYGON 5.655 0.67 5.19 0.67 5.19 0.32 5.25 0.32 5.25 0.61 5.595 0.61 5.595 0.32 5.655 0.32 ;
      RECT 4.985 0.32 5.045 1.345 ;
      RECT 4.295 2.385 4.74 2.445 ;
      POLYGON 4.735 1.13 4.465 1.13 4.465 0.25 4.455 0.25 4.455 0.23 4.44 0.23 4.44 0.17 4.455 0.17 4.455 0.13 4.515 0.13 4.515 0.17 4.525 0.17 4.525 1.07 4.735 1.07 ;
      RECT 4.645 0.135 4.705 0.995 ;
      POLYGON 4.395 1.51 4.135 1.51 4.135 0.83 3.6 0.83 3.6 0.245 3.66 0.245 3.66 0.77 4.135 0.77 4.135 0.32 4.195 0.32 4.195 1.45 4.395 1.45 ;
      POLYGON 4.205 3.17 4.145 3.17 4.145 2.78 3.345 2.78 3.345 2.72 4.145 2.72 4.145 2 4.205 2 ;
      POLYGON 4 2.93 3.27 2.93 3.27 3.17 3.21 3.17 3.21 2 3.27 2 3.27 2.87 4 2.87 ;
      RECT 3.71 1.24 3.99 1.525 ;
      RECT 3.415 0.32 3.475 1.455 ;
      POLYGON 3.27 1.52 2.935 1.52 2.935 1.46 3.21 1.46 3.21 0.32 3.27 0.32 ;
      RECT 2.675 0.6 2.735 1.29 ;
      POLYGON 2.445 0.83 2.385 0.83 2.385 1.485 2.325 1.485 2.325 0.32 2.385 0.32 2.385 0.77 2.445 0.77 ;
      POLYGON 2.385 3.085 2.325 3.085 2.325 2.74 1.855 2.74 1.855 2.68 2.325 2.68 2.325 2.185 2.385 2.185 ;
      POLYGON 2.265 1.19 2.18 1.19 2.18 1.485 2.12 1.485 2.12 1.13 2.205 1.13 2.205 0.585 1.51 0.585 1.51 1.27 1.63 1.27 1.63 1.485 1.295 1.485 1.295 1.27 1.45 1.27 1.45 0.585 1.115 0.585 1.115 0.595 1.085 0.595 1.085 1.14 1.115 1.14 1.115 1.2 0.995 1.2 0.995 1.14 1.025 1.14 1.025 0.595 0.995 0.595 0.995 0.535 1.025 0.535 1.025 0.525 1.675 0.525 1.675 0.32 1.735 0.32 1.735 0.525 2.12 0.525 2.12 0.32 2.18 0.32 2.18 0.525 2.265 0.525 ;
      POLYGON 2.115 0.705 2.075 0.705 2.075 0.75 2.06 0.75 2.06 1.18 2 1.18 2 0.705 1.995 0.705 1.995 0.645 2.115 0.645 ;
      POLYGON 1.975 0.465 1.915 0.465 1.915 0.255 1.53 0.255 1.53 0.465 1.47 0.465 1.47 0.195 1.975 0.195 ;
      POLYGON 1.915 0.705 1.885 0.705 1.885 1.185 1.725 1.185 1.725 1.2 1.605 1.2 1.605 1.14 1.635 1.14 1.635 1.125 1.825 1.125 1.825 0.705 1.795 0.705 1.795 0.645 1.915 0.645 ;
      POLYGON 1.87 2.535 1.745 2.535 1.745 2.875 1.87 2.875 1.87 3.085 1.81 3.085 1.81 2.935 1.685 2.935 1.685 2.475 1.81 2.475 1.81 2.24 1.39 2.24 1.39 2.2 1.255 2.2 1.255 1.955 0.665 1.955 0.665 3.115 0.605 3.115 0.605 1.895 1.315 1.895 1.315 2.14 1.45 2.14 1.45 2.18 1.87 2.18 ;
      POLYGON 1.315 3.115 1.255 3.115 1.255 2.605 0.975 2.605 0.975 2.545 1.255 2.545 1.255 2.28 1.315 2.28 ;
      POLYGON 0.905 3.115 0.845 3.115 0.845 2.115 0.75 2.115 0.75 2.055 0.905 2.055 ;
      POLYGON 0.84 1.485 0.43 1.485 0.43 1.56 0.37 1.56 0.37 1.425 0.78 1.425 0.78 0.32 0.84 0.32 ;
      RECT 0.61 0.135 0.67 1.305 ;
      POLYGON 0.55 0.985 0.51 0.985 0.51 1.265 0.45 1.265 0.45 0.32 0.51 0.32 0.51 0.865 0.55 0.865 ;
      POLYGON 0.46 3.115 0.4 3.115 0.4 1.965 0.34 1.965 0.34 1.905 0.46 1.905 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END SRDFFSRQX1

MACRO SRDFFSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SRDFFSRX1 0 0 ;
  SIZE 6.2 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 1.77 5.93 1.77 5.93 2.46 5.87 2.46 5.87 1.77 5.25 1.77 5.25 2.48 5.19 2.48 5.19 1.77 2.18 1.77 2.18 2.4 2.12 2.4 2.12 1.77 1.53 1.77 1.53 2.08 1.47 2.08 1.47 1.77 -0.005 1.77 -0.005 1.65 0.245 1.65 0.245 1.05 0.305 1.05 0.305 1.65 1.09 1.65 1.09 1.27 1.15 1.27 1.15 1.65 1.88 1.65 1.88 1.27 1.94 1.27 1.94 1.65 5.43 1.65 5.43 1.13 5.49 1.13 5.49 1.65 5.945 1.65 5.945 1.13 6.005 1.13 6.005 1.65 6.2 1.65 ;
    END
  END VDD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.26 2.585 2.255 2.585 2.255 2.605 2.02 2.605 2.02 2.465 2.255 2.465 2.255 2.525 2.26 2.525 ;
    END
  END SE
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0516 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.5925925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 23.37962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.37 0.925 1.29 0.925 1.29 1.14 1.32 1.14 1.32 1.2 1.2 1.2 1.2 1.14 1.23 1.14 1.23 0.925 1.225 0.925 1.225 0.72 1.37 0.72 ;
    END
  END SN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.895 2.61 3.415 2.61 3.415 2 3.545 2 3.545 1.89 3.795 1.89 3.795 2 3.895 2 ;
    END
  END ExtVDD
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.925926 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.385 0.905 0.375 0.905 0.375 0.935 0.245 0.935 0.245 0.755 0.375 0.755 0.375 0.845 0.385 0.845 ;
    END
  END RN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.673225 LAYER Metal1 ;
    ANTENNADIFFAREA 4.2416 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3015 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.81666675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 142.4179105 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.77 2.82 5.725 2.82 5.725 3.135 5.665 3.135 5.665 2.82 5.62 2.82 5.62 2.68 5.665 2.68 5.665 2.07 5.725 2.07 5.725 2.68 5.77 2.68 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.673225 LAYER Metal1 ;
    ANTENNADIFFAREA 4.271325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.3015 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.81666675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 142.4179105 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.045 3.13 4.985 3.13 4.985 2.855 4.805 2.855 4.805 2.67 4.985 2.67 4.985 2.09 5.045 2.09 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.574074 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.415 2.66 1.61 2.82 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.95 2.8 2.245 2.87 ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 3.48 0 3.48 0 3.36 1.05 3.36 1.05 2.97 1.11 2.97 1.11 3.36 1.5 3.36 1.5 2.94 1.56 2.94 1.56 3.36 2.12 3.36 2.12 2.94 2.18 2.94 2.18 3.36 3.415 3.36 3.415 3.025 3.475 3.025 3.475 3.36 3.835 3.36 3.835 3.025 3.895 3.025 3.895 3.36 5.19 3.36 5.19 2.87 5.25 2.87 5.25 3.36 5.87 3.36 5.87 2.875 5.93 2.875 5.93 3.36 6.2 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6.2 0.06 6.065 0.06 6.065 0.465 6.005 0.465 6.005 0.06 3.99 0.06 3.99 0.465 3.93 0.465 3.93 0.06 1.15 0.06 1.15 0.32 1.325 0.32 1.325 0.465 1.09 0.465 1.09 0.06 0.305 0.06 0.305 0.465 0.245 0.465 0.245 0.06 0 0.06 0 -0.06 6.2 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.58333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.77 1.525 4.455 1.525 4.455 1.37 4.31 1.37 4.31 0.41 4.37 0.41 4.37 1.31 4.77 1.31 ;
    END
  END RT
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.20370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.975 2.715 1.18 2.845 ;
    END
  END CK
  OBS
    LAYER Metal1 ;
      POLYGON 5.86 0.465 5.8 0.465 5.8 0.26 5.45 0.26 5.45 0.465 5.39 0.465 5.39 0.2 5.86 0.2 ;
      POLYGON 5.8 1.345 5.74 1.345 5.74 1.015 5.25 1.015 5.25 1.345 5.19 1.345 5.19 0.955 5.8 0.955 ;
      POLYGON 5.655 0.67 5.19 0.67 5.19 0.32 5.25 0.32 5.25 0.61 5.595 0.61 5.595 0.32 5.655 0.32 ;
      POLYGON 5.485 3.07 5.425 3.07 5.425 2.71 5.13 2.71 5.13 2.65 5.425 2.65 5.425 2.175 5.485 2.175 ;
      RECT 4.985 0.32 5.045 1.345 ;
      RECT 4.295 2.385 4.74 2.445 ;
      POLYGON 4.735 1.13 4.465 1.13 4.465 0.25 4.455 0.25 4.455 0.23 4.44 0.23 4.44 0.17 4.455 0.17 4.455 0.13 4.515 0.13 4.515 0.17 4.525 0.17 4.525 1.07 4.735 1.07 ;
      RECT 4.645 0.135 4.705 0.995 ;
      POLYGON 4.395 1.51 4.135 1.51 4.135 0.83 3.6 0.83 3.6 0.245 3.66 0.245 3.66 0.77 4.135 0.77 4.135 0.32 4.195 0.32 4.195 1.45 4.395 1.45 ;
      POLYGON 4.205 3.17 4.145 3.17 4.145 2.78 3.345 2.78 3.345 2.72 4.145 2.72 4.145 2 4.205 2 ;
      POLYGON 4 2.93 3.27 2.93 3.27 3.17 3.21 3.17 3.21 2 3.27 2 3.27 2.87 4 2.87 ;
      RECT 3.71 1.24 3.99 1.525 ;
      RECT 3.415 0.32 3.475 1.455 ;
      POLYGON 3.27 1.52 2.935 1.52 2.935 1.46 3.21 1.46 3.21 0.32 3.27 0.32 ;
      RECT 2.675 0.6 2.735 1.29 ;
      POLYGON 2.445 0.83 2.385 0.83 2.385 1.485 2.325 1.485 2.325 0.32 2.385 0.32 2.385 0.77 2.445 0.77 ;
      POLYGON 2.385 3.085 2.325 3.085 2.325 2.74 1.855 2.74 1.855 2.68 2.325 2.68 2.325 2.185 2.385 2.185 ;
      POLYGON 2.265 1.19 2.18 1.19 2.18 1.485 2.12 1.485 2.12 1.13 2.205 1.13 2.205 0.585 1.51 0.585 1.51 1.27 1.63 1.27 1.63 1.485 1.295 1.485 1.295 1.27 1.45 1.27 1.45 0.585 1.115 0.585 1.115 0.595 1.085 0.595 1.085 1.14 1.115 1.14 1.115 1.2 0.995 1.2 0.995 1.14 1.025 1.14 1.025 0.595 0.995 0.595 0.995 0.535 1.025 0.535 1.025 0.525 1.675 0.525 1.675 0.32 1.735 0.32 1.735 0.525 2.12 0.525 2.12 0.32 2.18 0.32 2.18 0.525 2.265 0.525 ;
      POLYGON 2.115 0.705 2.075 0.705 2.075 0.75 2.06 0.75 2.06 1.18 2 1.18 2 0.705 1.995 0.705 1.995 0.645 2.115 0.645 ;
      POLYGON 1.975 0.465 1.915 0.465 1.915 0.255 1.53 0.255 1.53 0.465 1.47 0.465 1.47 0.195 1.975 0.195 ;
      POLYGON 1.915 0.705 1.885 0.705 1.885 1.185 1.725 1.185 1.725 1.2 1.605 1.2 1.605 1.14 1.635 1.14 1.635 1.125 1.825 1.125 1.825 0.705 1.795 0.705 1.795 0.645 1.915 0.645 ;
      POLYGON 1.87 2.535 1.745 2.535 1.745 2.875 1.87 2.875 1.87 3.085 1.81 3.085 1.81 2.935 1.685 2.935 1.685 2.475 1.81 2.475 1.81 2.24 1.39 2.24 1.39 2.2 1.255 2.2 1.255 1.93 0.665 1.93 0.665 3.115 0.605 3.115 0.605 1.87 1.315 1.87 1.315 2.14 1.45 2.14 1.45 2.18 1.87 2.18 ;
      POLYGON 1.315 3.115 1.255 3.115 1.255 2.625 0.97 2.625 0.97 2.565 1.255 2.565 1.255 2.28 1.315 2.28 ;
      POLYGON 0.905 3.115 0.845 3.115 0.845 2.105 0.77 2.105 0.77 2.045 0.905 2.045 ;
      POLYGON 0.84 1.485 0.43 1.485 0.43 1.56 0.37 1.56 0.37 1.425 0.78 1.425 0.78 0.32 0.84 0.32 ;
      RECT 0.61 0.135 0.67 1.305 ;
      POLYGON 0.55 0.985 0.51 0.985 0.51 1.265 0.45 1.265 0.45 0.32 0.51 0.32 0.51 0.865 0.55 0.865 ;
      POLYGON 0.46 3.115 0.4 3.115 0.4 1.965 0.34 1.965 0.34 1.905 0.46 1.905 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END SRDFFSRX1

MACRO SRDFFSX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SRDFFSX1 0 0 ;
  SIZE 6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 1.77 5.73 1.77 5.73 2.46 5.67 2.46 5.67 1.77 5.05 1.77 5.05 2.48 4.99 2.48 4.99 1.77 1.98 1.77 1.98 2.4 1.92 2.4 1.92 1.77 1.33 1.77 1.33 2.08 1.27 2.08 1.27 1.77 -0.005 1.77 -0.005 1.65 0.89 1.65 0.89 1.27 0.95 1.27 0.95 1.65 1.575 1.65 1.575 1.27 1.635 1.27 1.635 1.65 5.23 1.65 5.23 1.13 5.29 1.13 5.29 1.65 5.64 1.65 5.64 1.13 5.7 1.13 5.7 1.65 6 1.65 ;
    END
  END VDD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.06 2.585 2.055 2.585 2.055 2.605 1.82 2.605 1.82 2.465 2.055 2.465 2.055 2.525 2.06 2.525 ;
    END
  END SE
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0516 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.5925925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 23.37962975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.17 0.945 1.09 0.945 1.09 1.14 1.12 1.14 1.12 1.2 1 1.2 1 1.14 1.03 1.14 1.03 0.945 1.025 0.945 1.025 0.72 1.17 0.72 ;
    END
  END SN
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.695 2.61 3.215 2.61 3.215 2 3.345 2 3.345 1.89 3.595 1.89 3.595 2 3.695 2 ;
    END
  END ExtVDD
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.257875 LAYER Metal1 ;
    ANTENNADIFFAREA 3.9742 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2691 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.53874025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 145.039019 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.57 2.83 5.525 2.83 5.525 3.135 5.465 3.135 5.465 2.83 5.405 2.83 5.405 2.67 5.465 2.67 5.465 2.07 5.525 2.07 5.525 2.67 5.57 2.67 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.257875 LAYER Metal1 ;
    ANTENNADIFFAREA 3.9742 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2691 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.53874025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 145.039019 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.845 3.13 4.785 3.13 4.785 2.82 4.62 2.82 4.62 2.685 4.785 2.685 4.785 2.09 4.845 2.09 ;
    END
  END QN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.5555555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.78 2.745 0.98 2.845 ;
    END
  END CK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 2.66 1.41 2.79 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.75 2.8 2.045 2.87 ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 3.48 0 3.48 0 3.36 0.85 3.36 0.85 2.97 0.91 2.97 0.91 3.36 1.3 3.36 1.3 2.94 1.36 2.94 1.36 3.36 1.92 3.36 1.92 2.94 1.98 2.94 1.98 3.36 3.215 3.36 3.215 3.025 3.275 3.025 3.275 3.36 3.635 3.36 3.635 3.025 3.695 3.025 3.695 3.36 4.99 3.36 4.99 2.87 5.05 2.87 5.05 3.36 5.67 3.36 5.67 2.875 5.73 2.875 5.73 3.36 6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6 0.06 5.265 0.06 5.265 0.35 5.26 0.35 5.26 0.465 5.2 0.465 5.2 0.32 5.205 0.32 5.205 0.06 3.79 0.06 3.79 0.465 3.73 0.465 3.73 0.06 0.95 0.06 0.95 0.32 1.185 0.32 1.185 0.44 1.125 0.44 1.125 0.465 0.89 0.465 0.89 0.06 0 0.06 0 -0.06 6 -0.06 ;
    END
  END VSS
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.10185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.41 1.525 4.255 1.525 4.255 1.37 4.11 1.37 4.11 0.41 4.17 0.41 4.17 1.31 4.41 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.495 1.345 5.435 1.345 5.435 1.015 5.05 1.015 5.05 1.345 4.99 1.345 4.99 0.955 5.495 0.955 ;
      POLYGON 5.285 3.07 5.225 3.07 5.225 2.71 4.93 2.71 4.93 2.65 5.225 2.65 5.225 2.175 5.285 2.175 ;
      RECT 4.785 0.32 4.845 1.345 ;
      RECT 4.095 2.385 4.54 2.445 ;
      POLYGON 4.535 1.13 4.265 1.13 4.265 0.25 4.255 0.25 4.255 0.23 4.24 0.23 4.24 0.17 4.255 0.17 4.255 0.13 4.315 0.13 4.315 0.17 4.325 0.17 4.325 1.07 4.535 1.07 ;
      RECT 4.445 0.135 4.505 0.995 ;
      POLYGON 4.195 1.51 3.935 1.51 3.935 0.83 3.4 0.83 3.4 0.245 3.46 0.245 3.46 0.77 3.935 0.77 3.935 0.32 3.995 0.32 3.995 1.45 4.195 1.45 ;
      POLYGON 4.005 3.17 3.945 3.17 3.945 2.78 3.145 2.78 3.145 2.72 3.945 2.72 3.945 2 4.005 2 ;
      POLYGON 3.8 2.93 3.07 2.93 3.07 3.17 3.01 3.17 3.01 2 3.07 2 3.07 2.87 3.8 2.87 ;
      RECT 3.51 1.24 3.79 1.525 ;
      RECT 3.215 0.32 3.275 1.455 ;
      POLYGON 3.07 1.52 2.735 1.52 2.735 1.46 3.01 1.46 3.01 0.32 3.07 0.32 ;
      RECT 2.475 0.6 2.535 1.29 ;
      POLYGON 2.245 0.83 2.185 0.83 2.185 1.485 2.125 1.485 2.125 0.32 2.185 0.32 2.185 0.77 2.245 0.77 ;
      POLYGON 2.185 3.085 2.125 3.085 2.125 2.74 1.655 2.74 1.655 2.68 2.125 2.68 2.125 2.185 2.185 2.185 ;
      POLYGON 1.98 1.485 1.92 1.485 1.92 0.585 1.31 0.585 1.31 1.27 1.43 1.27 1.43 1.485 1.095 1.485 1.095 1.27 1.25 1.27 1.25 0.585 0.915 0.585 0.915 0.595 0.885 0.595 0.885 1.14 0.915 1.14 0.915 1.2 0.795 1.2 0.795 1.14 0.825 1.14 0.825 0.595 0.795 0.595 0.795 0.535 0.825 0.535 0.825 0.525 1.475 0.525 1.475 0.32 1.535 0.32 1.535 0.525 1.92 0.525 1.92 0.32 1.98 0.32 ;
      POLYGON 1.715 0.705 1.685 0.705 1.685 1.185 1.525 1.185 1.525 1.2 1.405 1.2 1.405 1.14 1.435 1.14 1.435 1.125 1.625 1.125 1.625 0.705 1.595 0.705 1.595 0.645 1.715 0.645 ;
      POLYGON 1.67 2.535 1.545 2.535 1.545 2.875 1.67 2.875 1.67 3.085 1.61 3.085 1.61 2.935 1.485 2.935 1.485 2.475 1.61 2.475 1.61 2.24 1.19 2.24 1.19 2.2 1.055 2.2 1.055 1.93 0.465 1.93 0.465 3.115 0.405 3.115 0.405 1.87 1.115 1.87 1.115 2.14 1.25 2.14 1.25 2.18 1.67 2.18 ;
      POLYGON 1.115 3.115 1.055 3.115 1.055 2.64 0.775 2.64 0.775 2.58 1.055 2.58 1.055 2.28 1.115 2.28 ;
      POLYGON 0.705 3.115 0.645 3.115 0.645 2.105 0.535 2.105 0.535 2.045 0.705 2.045 ;
      POLYGON 0.64 1.485 0.23 1.485 0.23 1.56 0.17 1.56 0.17 1.425 0.58 1.425 0.58 0.32 0.64 0.32 ;
      RECT 0.41 0.135 0.47 1.305 ;
      POLYGON 0.26 3.115 0.2 3.115 0.2 1.965 0.14 1.965 0.14 1.905 0.26 1.905 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END SRDFFSX1

MACRO SRDFFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SRDFFX1 0 0 ;
  SIZE 6 BY 3.42 ;
  SYMMETRY X Y ;
  SITE CoreSiteDouble ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 1.77 5.73 1.77 5.73 2.46 5.67 2.46 5.67 1.77 5.05 1.77 5.05 2.48 4.99 2.48 4.99 1.77 1.98 1.77 1.98 2.4 1.92 2.4 1.92 1.77 1.33 1.77 1.33 2.08 1.27 2.08 1.27 1.77 -0.005 1.77 -0.005 1.65 0.89 1.65 0.89 1.27 0.95 1.27 0.95 1.65 5.23 1.65 5.23 1.13 5.29 1.13 5.29 1.65 6 1.65 ;
    END
  END VDD
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.06 2.585 2.055 2.585 2.055 2.605 1.82 2.605 1.82 2.465 2.055 2.465 2.055 2.525 2.06 2.525 ;
    END
  END SE
  PIN ExtVDD
    DIRECTION INOUT ;
    USE POWER ;
    NETEXPR "ExtVDD ExtVDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.695 2.61 3.215 2.61 3.215 2 3.345 2 3.345 1.89 3.595 1.89 3.595 2 3.695 2 ;
    END
  END ExtVDD
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.06 LAYER Metal1 ;
    ANTENNADIFFAREA 3.822325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2691 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.80341875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 139.7324415 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.565 2.625 5.525 2.625 5.525 3.135 5.465 3.135 5.465 2.625 5.375 2.625 5.375 2.495 5.465 2.495 5.465 2.07 5.525 2.07 5.525 2.495 5.565 2.495 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.06 LAYER Metal1 ;
    ANTENNADIFFAREA 3.822325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2691 LAYER Metal1 ;
      ANTENNAMAXAREACAR 18.80341875 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 139.7324415 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.845 3.13 4.785 3.13 4.785 2.83 4.62 2.83 4.62 2.67 4.785 2.67 4.785 2.09 4.845 2.09 ;
    END
  END QN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.215 2.66 1.41 2.79 ;
    END
  END D
  PIN SI
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.75 2.8 2.045 2.87 ;
    END
  END SI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6 3.48 0 3.48 0 3.36 0.85 3.36 0.85 2.97 0.91 2.97 0.91 3.36 1.3 3.36 1.3 2.94 1.36 2.94 1.36 3.36 1.92 3.36 1.92 2.94 1.98 2.94 1.98 3.36 3.215 3.36 3.215 3.025 3.275 3.025 3.275 3.36 3.635 3.36 3.635 3.025 3.695 3.025 3.695 3.36 4.99 3.36 4.99 2.87 5.05 2.87 5.05 3.36 5.67 3.36 5.67 2.875 5.73 2.875 5.73 3.36 6 3.36 ;
    END
    PORT
      LAYER Metal1 ;
        POLYGON 6 0.06 5.155 0.06 5.155 0.465 5.095 0.465 5.095 0.06 3.79 0.06 3.79 0.465 3.73 0.465 3.73 0.06 0.95 0.06 0.95 0.465 0.89 0.465 0.89 0.06 0 0.06 0 -0.06 6 -0.06 ;
    END
  END VSS
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.64814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.775 2.745 0.98 2.845 ;
    END
  END CK
  PIN RT
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 14.7685185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.59 1.525 4.255 1.525 4.255 1.37 4.11 1.37 4.11 0.41 4.17 0.41 4.17 1.31 4.59 1.31 ;
    END
  END RT
  OBS
    LAYER Metal1 ;
      POLYGON 5.495 1.345 5.435 1.345 5.435 1.015 5.05 1.015 5.05 1.345 4.99 1.345 4.99 0.955 5.495 0.955 ;
      POLYGON 5.285 3.07 5.225 3.07 5.225 2.71 4.93 2.71 4.93 2.65 5.225 2.65 5.225 2.175 5.285 2.175 ;
      RECT 4.785 0.32 4.845 1.345 ;
      RECT 4.095 2.385 4.54 2.445 ;
      POLYGON 4.535 1.07 4.265 1.07 4.265 0.25 4.255 0.25 4.255 0.23 4.24 0.23 4.24 0.17 4.255 0.17 4.255 0.13 4.315 0.13 4.315 0.17 4.325 0.17 4.325 1.01 4.535 1.01 ;
      POLYGON 4.195 1.51 3.935 1.51 3.935 0.83 3.4 0.83 3.4 0.245 3.46 0.245 3.46 0.77 3.935 0.77 3.935 0.32 3.995 0.32 3.995 1.45 4.195 1.45 ;
      POLYGON 4.005 3.17 3.945 3.17 3.945 2.78 3.145 2.78 3.145 2.72 3.945 2.72 3.945 2 4.005 2 ;
      POLYGON 3.8 2.93 3.07 2.93 3.07 3.17 3.01 3.17 3.01 2 3.07 2 3.07 2.87 3.8 2.87 ;
      RECT 3.51 1.24 3.79 1.525 ;
      RECT 3.215 0.32 3.275 1.455 ;
      POLYGON 3.07 1.52 2.735 1.52 2.735 1.46 3.01 1.46 3.01 0.32 3.07 0.32 ;
      RECT 2.475 0.6 2.535 1.29 ;
      POLYGON 2.245 0.83 2.185 0.83 2.185 1.485 2.125 1.485 2.125 0.32 2.185 0.32 2.185 0.77 2.245 0.77 ;
      POLYGON 2.185 3.085 2.125 3.085 2.125 2.74 1.655 2.74 1.655 2.68 2.125 2.68 2.125 2.185 2.185 2.185 ;
      POLYGON 1.98 1.485 1.92 1.485 1.92 0.585 1.155 0.585 1.155 1.485 1.095 1.485 1.095 0.585 0.915 0.585 0.915 0.595 0.885 0.595 0.885 1.14 0.915 1.14 0.915 1.2 0.795 1.2 0.795 1.14 0.825 1.14 0.825 0.595 0.795 0.595 0.795 0.535 0.825 0.535 0.825 0.525 1.095 0.525 1.095 0.32 1.155 0.32 1.155 0.525 1.92 0.525 1.92 0.32 1.98 0.32 ;
      POLYGON 1.67 2.535 1.545 2.535 1.545 2.875 1.67 2.875 1.67 3.085 1.61 3.085 1.61 2.935 1.485 2.935 1.485 2.475 1.61 2.475 1.61 2.24 1.19 2.24 1.19 2.2 1.055 2.2 1.055 1.93 0.465 1.93 0.465 3.115 0.405 3.115 0.405 1.87 1.115 1.87 1.115 2.14 1.25 2.14 1.25 2.18 1.67 2.18 ;
      POLYGON 1.115 3.115 1.055 3.115 1.055 2.64 0.775 2.64 0.775 2.58 1.055 2.58 1.055 2.28 1.115 2.28 ;
      POLYGON 0.705 3.115 0.645 3.115 0.645 2.105 0.57 2.105 0.57 2.045 0.705 2.045 ;
      POLYGON 0.64 1.485 0.23 1.485 0.23 1.56 0.17 1.56 0.17 1.425 0.58 1.425 0.58 0.32 0.64 0.32 ;
      RECT 0.41 0.135 0.47 1.305 ;
      POLYGON 0.26 3.115 0.2 3.115 0.2 1.965 0.14 1.965 0.14 1.905 0.26 1.905 ;
  END
  PROPERTY oaTaper "virtuosoDefaultTaper" ;
END SRDFFX1

MACRO TBUFX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX1 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.03515 LAYER Metal1 ;
    ANTENNADIFFAREA 1.120875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXAREACAR 22.7755775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 173.59735975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.965 1.3 1.87 1.3 1.87 0.91 1.905 0.91 1.905 0.555 1.735 0.555 1.735 0.435 1.965 0.435 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 18.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.43 0.345 1.29 0.345 1.29 0.37 0.78 0.37 0.78 0.665 0.88 0.665 0.88 1.065 0.765 1.065 0.765 1.085 0.635 1.085 0.635 1.065 0.43 1.065 0.43 1.005 0.82 1.005 0.82 0.725 0.72 0.725 0.72 0.31 1.23 0.31 1.23 0.285 1.43 0.285 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.54629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.72 0.905 0.33 0.905 0.33 0.945 0.25 0.945 0.25 0.825 0.46 0.825 0.46 0.6 0.54 0.6 0.54 0.825 0.72 0.825 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.11 1.65 0.11 1.24 0.17 1.24 0.17 1.65 0.53 1.65 0.53 1.54 0.65 1.54 0.65 1.65 1.655 1.65 1.655 0.975 1.715 0.975 1.715 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.59 0.06 1.59 0.42 1.53 0.42 1.53 0.06 1.13 0.06 1.13 0.17 1.01 0.17 1.01 0.06 0.62 0.06 0.62 0.5 0.56 0.5 0.56 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.77 0.875 1.555 0.875 1.555 1.405 0.325 1.405 0.325 1.225 0.27 1.225 0.27 1.14 0.09 1.14 0.09 0.56 0.175 0.56 0.175 0.5 0.235 0.5 0.235 0.62 0.15 0.62 0.15 1.08 0.33 1.08 0.33 1.165 0.385 1.165 0.385 1.345 1.495 1.345 1.495 0.815 1.71 0.815 1.71 0.74 1.77 0.74 ;
      POLYGON 1.61 0.715 1.395 0.715 1.395 0.86 1.26 0.86 1.26 1 1.14 1 1.14 0.94 1.2 0.94 1.2 0.8 1.335 0.8 1.335 0.53 1.245 0.53 1.245 0.47 1.395 0.47 1.395 0.655 1.61 0.655 ;
      POLYGON 1.235 0.7 1.04 0.7 1.04 1.245 0.765 1.245 0.765 1.185 0.98 1.185 0.98 0.565 0.88 0.565 0.88 0.505 1.04 0.505 1.04 0.64 1.235 0.64 ;
  END
END TBUFX1

MACRO TBUFX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX12 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5223 LAYER Metal1 ;
    ANTENNADIFFAREA 4.574 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.4383 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.0362765 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 62.587269 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.325 1.405 6.265 1.405 6.265 0.92 5.915 0.92 5.915 1.405 5.855 1.405 5.855 0.92 5.505 0.92 5.505 1.405 5.445 1.405 5.445 0.92 5.095 0.92 5.095 1.405 5.035 1.405 5.035 0.92 4.685 0.92 4.685 1.405 4.625 1.405 4.625 0.92 4.32 0.92 4.32 1.08 4.275 1.08 4.275 1.405 4.215 1.405 4.215 1.02 4.26 1.02 4.26 0.555 4.1 0.555 4.1 0.415 4.16 0.415 4.16 0.495 4.32 0.495 4.32 0.79 4.34 0.79 4.34 0.86 4.625 0.86 4.625 0.555 4.51 0.555 4.51 0.415 4.57 0.415 4.57 0.495 4.92 0.495 4.92 0.415 4.98 0.415 4.98 0.555 4.685 0.555 4.685 0.86 5.855 0.86 5.855 0.555 5.33 0.555 5.33 0.415 5.39 0.415 5.39 0.495 5.74 0.495 5.74 0.415 5.8 0.415 5.8 0.495 6.15 0.495 6.15 0.415 6.21 0.415 6.21 0.555 5.915 0.555 5.915 0.86 6.325 0.86 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1746 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.694158 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.78 0.865 2.36 0.865 2.36 0.705 2.065 0.705 2.065 0.35 1.72 0.35 1.72 0.675 1.28 0.675 1.28 0.355 0.96 0.355 0.96 0.865 0.765 0.865 0.765 0.895 0.635 0.895 0.635 0.865 0.54 0.865 0.54 0.805 0.9 0.805 0.9 0.295 1.34 0.295 1.34 0.615 1.66 0.615 1.66 0.29 2.125 0.29 2.125 0.645 2.42 0.645 2.42 0.805 3.72 0.805 3.72 0.745 3.78 0.745 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.05 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.11655 LAYER Metal1 ;
      ANTENNAMAXAREACAR 0.4290005 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.26383525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 0.705 0.44 0.705 0.44 0.78 0.36 0.78 0.36 0.625 0.72 0.625 0.72 0.585 0.8 0.585 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 1.77 0 1.77 0 1.65 0.435 1.65 0.435 1.315 0.555 1.315 0.555 1.375 0.495 1.375 0.495 1.65 0.935 1.65 0.935 1.51 0.995 1.51 0.995 1.65 1.51 1.65 1.51 1.51 1.57 1.51 1.57 1.65 1.91 1.65 1.91 1.51 1.97 1.51 1.97 1.65 2.365 1.65 2.365 1.51 2.425 1.51 2.425 1.65 3.125 1.65 3.125 1.285 3.245 1.285 3.245 1.345 3.185 1.345 3.185 1.65 3.905 1.65 3.905 1.285 3.965 1.285 3.965 1.65 4.42 1.65 4.42 1.02 4.48 1.02 4.48 1.65 4.83 1.65 4.83 1.02 4.89 1.02 4.89 1.65 5.24 1.65 5.24 1.02 5.3 1.02 5.3 1.65 5.65 1.65 5.65 1.02 5.71 1.02 5.71 1.65 6.06 1.65 6.06 1.02 6.12 1.02 6.12 1.65 6.47 1.65 6.47 1.015 6.53 1.015 6.53 1.65 6.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 0.06 6.415 0.06 6.415 0.395 6.355 0.395 6.355 0.06 6.005 0.06 6.005 0.395 5.945 0.395 5.945 0.06 5.595 0.06 5.595 0.395 5.535 0.395 5.535 0.06 5.185 0.06 5.185 0.395 5.125 0.395 5.125 0.06 4.775 0.06 4.775 0.395 4.715 0.395 4.715 0.06 4.365 0.06 4.365 0.395 4.305 0.395 4.305 0.06 3.955 0.06 3.955 0.395 3.895 0.395 3.895 0.06 3.515 0.06 3.515 0.305 3.575 0.305 3.575 0.365 3.455 0.365 3.455 0.06 3.105 0.06 3.105 0.305 3.165 0.305 3.165 0.365 3.045 0.365 3.045 0.06 2.695 0.06 2.695 0.305 2.755 0.305 2.755 0.365 2.635 0.365 2.635 0.06 2.345 0.06 2.345 0.44 2.225 0.44 2.225 0.38 2.285 0.38 2.285 0.06 1.56 0.06 1.56 0.44 1.44 0.44 1.44 0.38 1.5 0.38 1.5 0.06 0.495 0.06 0.495 0.47 0.435 0.47 0.435 0.06 0 0.06 0 -0.06 6.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.16 0.92 4.1 0.92 4.1 1.185 3.805 1.185 3.805 1.395 3.425 1.395 3.425 1.185 2.145 1.185 2.145 1.055 0.67 1.055 0.67 0.995 1.06 0.995 1.06 0.455 1.18 0.455 1.18 0.515 1.12 0.515 1.12 0.995 1.905 0.995 1.905 0.51 1.82 0.51 1.82 0.45 1.965 0.45 1.965 0.995 2.205 0.995 2.205 1.125 3.485 1.125 3.485 1.335 3.745 1.335 3.745 1.125 4.04 1.125 4.04 0.86 4.16 0.86 ;
      POLYGON 3.995 0.695 3.94 0.695 3.94 1.025 3.645 1.025 3.645 1.235 3.585 1.235 3.585 1.025 2.785 1.025 2.785 0.965 3.88 0.965 3.88 0.635 3.69 0.635 3.69 0.525 2.46 0.525 2.46 0.35 2.52 0.35 2.52 0.465 2.87 0.465 2.87 0.35 2.93 0.35 2.93 0.465 3.28 0.465 3.28 0.345 3.34 0.345 3.34 0.465 3.69 0.465 3.69 0.345 3.75 0.345 3.75 0.575 3.995 0.575 ;
      RECT 2.71 0.625 3.51 0.705 ;
      POLYGON 2.83 1.37 2.71 1.37 2.71 1.345 0.655 1.345 0.655 1.215 0.26 1.215 0.26 1.335 0.2 1.335 0.2 0.49 0.26 0.49 0.26 1.155 0.715 1.155 0.715 1.285 2.77 1.285 2.77 1.31 2.83 1.31 ;
      POLYGON 1.805 0.855 1.3 0.855 1.3 0.895 1.22 0.895 1.22 0.775 1.805 0.775 ;
  END
END TBUFX12

MACRO TBUFX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX16 0 0 ;
  SIZE 9 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.6098 LAYER Metal1 ;
    ANTENNADIFFAREA 5.978575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.583875 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.895183 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 60.660244 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.545 1.42 8.485 1.42 8.485 1.09 8.135 1.09 8.135 1.42 8.075 1.42 8.075 1.09 7.725 1.09 7.725 1.42 7.665 1.42 7.665 1.09 7.315 1.09 7.315 1.42 7.255 1.42 7.255 1.09 6.905 1.09 6.905 1.42 6.845 1.42 6.845 1.09 6.495 1.09 6.495 1.42 6.435 1.42 6.435 1.09 6.085 1.09 6.085 1.42 6.025 1.42 6.025 1.09 5.72 1.09 5.72 1.125 5.675 1.125 5.675 1.42 5.615 1.42 5.615 1.065 5.66 1.065 5.66 0.51 5.5 0.51 5.5 0.37 5.56 0.37 5.56 0.45 5.72 0.45 5.72 0.79 5.74 0.79 5.74 1.03 6.025 1.03 6.025 0.51 5.91 0.51 5.91 0.37 5.97 0.37 5.97 0.45 6.32 0.45 6.32 0.37 6.38 0.37 6.38 0.51 6.085 0.51 6.085 1.03 7.14 1.03 7.14 0.51 6.73 0.51 6.73 0.37 6.79 0.37 6.79 0.45 7.14 0.45 7.14 0.37 7.2 0.37 7.2 1.03 8.37 1.03 8.37 0.51 7.55 0.51 7.55 0.37 7.61 0.37 7.61 0.45 7.96 0.45 7.96 0.37 8.02 0.37 8.02 0.45 8.37 0.45 8.37 0.37 8.43 0.37 8.43 1.03 8.545 1.03 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.23175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.8478965 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.18 0.695 4.92 0.695 4.92 0.67 3.06 0.67 3.06 0.51 3.02 0.51 3.02 0.47 2.625 0.47 2.625 0.735 2.4 0.735 2.4 0.845 2.34 0.845 2.34 0.735 2.245 0.735 2.245 0.47 1.865 0.47 1.865 0.705 1.655 0.705 1.655 0.83 1.595 0.83 1.595 0.705 1.425 0.705 1.425 0.47 1.095 0.47 1.095 0.815 1.165 0.815 1.165 0.895 1.095 0.895 1.095 0.99 0.705 0.99 0.705 0.93 0.515 0.93 0.515 0.87 0.765 0.87 0.765 0.93 1.035 0.93 1.035 0.41 1.485 0.41 1.485 0.645 1.805 0.645 1.805 0.41 2.305 0.41 2.305 0.675 2.565 0.675 2.565 0.41 3.08 0.41 3.08 0.45 3.12 0.45 3.12 0.61 4.98 0.61 4.98 0.635 5.18 0.635 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.11955 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.145125 LAYER Metal1 ;
      ANTENNAMAXAREACAR 0.8237725 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.235142 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.935 0.83 0.875 0.83 0.875 0.77 0.415 0.77 0.415 0.92 0.26 0.92 0.26 0.71 0.935 0.71 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 9 1.77 0 1.77 0 1.65 0.25 1.65 0.25 1.255 0.31 1.255 0.31 1.65 0.69 1.65 0.69 1.51 0.75 1.51 0.75 1.65 1.26 1.65 1.26 1.255 1.32 1.255 1.32 1.65 1.7 1.65 1.7 1.51 1.76 1.51 1.76 1.65 2.14 1.65 2.14 1.255 2.2 1.255 2.2 1.65 2.58 1.65 2.58 1.26 2.52 1.26 2.52 1.2 2.64 1.2 2.64 1.65 3.765 1.65 3.765 1.25 3.885 1.25 3.885 1.31 3.825 1.31 3.825 1.65 4.465 1.65 4.465 1.25 4.585 1.25 4.585 1.31 4.525 1.31 4.525 1.65 5.165 1.65 5.165 1.25 5.285 1.25 5.285 1.31 5.225 1.31 5.225 1.65 5.82 1.65 5.82 1.19 5.88 1.19 5.88 1.65 6.23 1.65 6.23 1.19 6.29 1.19 6.29 1.65 6.64 1.65 6.64 1.19 6.7 1.19 6.7 1.65 7.05 1.65 7.05 1.19 7.11 1.19 7.11 1.65 7.46 1.65 7.46 1.19 7.52 1.19 7.52 1.65 7.87 1.65 7.87 1.19 7.93 1.19 7.93 1.65 8.28 1.65 8.28 1.19 8.34 1.19 8.34 1.65 8.69 1.65 8.69 1.03 8.75 1.03 8.75 1.65 9 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 9 0.06 8.635 0.06 8.635 0.35 8.575 0.35 8.575 0.06 8.225 0.06 8.225 0.35 8.165 0.35 8.165 0.06 7.815 0.06 7.815 0.35 7.755 0.35 7.755 0.06 7.405 0.06 7.405 0.35 7.345 0.35 7.345 0.06 6.995 0.06 6.995 0.35 6.935 0.35 6.935 0.06 6.585 0.06 6.585 0.35 6.525 0.35 6.525 0.06 6.175 0.06 6.175 0.35 6.115 0.35 6.115 0.06 5.765 0.06 5.765 0.35 5.705 0.35 5.705 0.06 5.33 0.06 5.33 0.35 5.27 0.35 5.27 0.06 4.92 0.06 4.92 0.35 4.86 0.35 4.86 0.06 4.51 0.06 4.51 0.35 4.45 0.35 4.45 0.06 4.06 0.06 4.06 0.35 4 0.35 4 0.06 3.65 0.06 3.65 0.35 3.59 0.35 3.59 0.06 3.24 0.06 3.24 0.35 3.18 0.35 3.18 0.06 2.465 0.06 2.465 0.575 2.405 0.575 2.405 0.06 1.645 0.06 1.645 0.485 1.705 0.485 1.705 0.545 1.585 0.545 1.585 0.06 0.68 0.06 0.68 0.575 0.62 0.575 0.62 0.06 0 0.06 0 -0.06 9 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.56 0.965 5.515 0.965 5.515 1.15 5.065 1.15 5.065 1.31 4.685 1.31 4.685 1.15 4.365 1.15 4.365 1.31 3.985 1.31 3.985 1.15 3.665 1.15 3.665 1.31 2.74 1.31 2.74 1.1 2.405 1.1 2.405 1.21 2.345 1.21 2.345 1.15 1.995 1.15 1.995 1.21 1.935 1.21 1.935 1.15 1.525 1.15 1.525 1.375 1.465 1.375 1.465 1.15 0.985 1.15 0.985 1.21 0.925 1.21 0.925 1.15 0.515 1.15 0.515 1.375 0.455 1.375 0.455 1.15 0.1 1.15 0.1 0.55 0.25 0.55 0.25 0.49 0.31 0.49 0.31 0.61 0.16 0.61 0.16 1.09 1.265 1.09 1.265 0.63 1.205 0.63 1.205 0.57 1.325 0.57 1.325 1.09 2.085 1.09 2.085 0.63 1.965 0.63 1.965 0.57 2.145 0.57 2.145 1.09 2.345 1.09 2.345 1.04 2.8 1.04 2.8 1.25 3.605 1.25 3.605 1.09 4.045 1.09 4.045 1.25 4.305 1.25 4.305 1.09 4.745 1.09 4.745 1.25 5.005 1.25 5.005 1.09 5.455 1.09 5.455 0.905 5.5 0.905 5.5 0.845 5.56 0.845 ;
      POLYGON 5.4 0.695 5.34 0.695 5.34 0.99 4.905 0.99 4.905 1.15 4.845 1.15 4.845 0.99 4.205 0.99 4.205 1.15 4.145 1.15 4.145 0.99 3.505 0.99 3.505 1.15 3.445 1.15 3.445 0.93 5.28 0.93 5.28 0.51 3.385 0.51 3.385 0.23 3.445 0.23 3.445 0.45 3.795 0.45 3.795 0.315 3.855 0.315 3.855 0.45 4.205 0.45 4.205 0.315 4.265 0.315 4.265 0.45 4.655 0.45 4.655 0.315 4.715 0.315 4.715 0.45 5.065 0.45 5.065 0.315 5.125 0.315 5.125 0.45 5.34 0.45 5.34 0.635 5.4 0.635 ;
      POLYGON 4.82 0.83 3.02 0.83 3.02 0.99 2.9 0.99 2.9 0.67 2.725 0.67 2.725 0.57 2.845 0.57 2.845 0.61 2.96 0.61 2.96 0.77 4.82 0.77 ;
      POLYGON 1.985 0.99 1.425 0.99 1.425 0.87 1.485 0.87 1.485 0.93 1.865 0.93 1.865 0.805 1.985 0.805 ;
  END
END TBUFX16

MACRO TBUFX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX2 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.1075 LAYER Metal1 ;
    ANTENNADIFFAREA 1.267775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0747 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.8259705 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 112.5301205 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 1.28 1.86 1.28 1.86 0.49 1.835 0.49 1.835 0.37 1.94 0.37 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 16.75925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.52 0.75 1.46 0.75 1.46 1.2 0.705 1.2 0.705 0.895 0.635 0.895 0.635 0.865 0.555 0.865 0.555 0.805 0.695 0.805 0.695 0.815 0.765 0.815 0.765 1.14 1.4 1.14 1.4 0.69 1.52 0.69 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.765 0.705 0.405 0.705 0.405 0.745 0.29 0.745 0.29 0.705 0.235 0.705 0.235 0.625 0.765 0.625 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.16 1.65 0.16 1.045 0.22 1.045 0.22 1.65 0.565 1.65 0.565 1.54 0.685 1.54 0.685 1.65 1.6 1.65 1.6 1.54 1.72 1.54 1.72 1.65 2.07 1.65 2.07 0.9 2.13 0.9 2.13 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 2.1 0.06 2.1 0.35 2.04 0.35 2.04 0.06 1.6 0.06 1.6 0.34 1.66 0.34 1.66 0.4 1.54 0.4 1.54 0.06 1.22 0.06 1.22 0.43 1.16 0.43 1.16 0.06 0.685 0.06 0.685 0.525 0.625 0.525 0.625 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.94 1.445 1.82 1.445 1.82 1.44 0.365 1.44 0.365 0.945 0.075 0.945 0.075 0.465 0.215 0.465 0.215 0.405 0.275 0.405 0.275 0.525 0.135 0.525 0.135 0.885 0.425 0.885 0.425 1.38 1.88 1.38 1.88 1.385 1.94 1.385 ;
      POLYGON 1.68 0.65 1.62 0.65 1.62 0.59 1.3 0.59 1.3 1.04 1.18 1.04 1.18 0.98 1.24 0.98 1.24 0.53 1.365 0.53 1.365 0.335 1.425 0.335 1.425 0.53 1.68 0.53 ;
      POLYGON 1.14 0.68 0.925 0.68 0.925 0.98 0.985 0.98 0.985 1.04 0.865 1.04 0.865 0.43 0.925 0.43 0.925 0.62 1.14 0.62 ;
  END
END TBUFX2

MACRO TBUFX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX20 0 0 ;
  SIZE 10 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.182425 LAYER Metal1 ;
    ANTENNADIFFAREA 7.23835 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.7308 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.091441 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 54.53612475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 9.725 1.415 9.665 1.415 9.665 1.085 9.315 1.085 9.315 1.415 9.255 1.415 9.255 1.085 8.905 1.085 8.905 1.415 8.845 1.415 8.845 1.085 8.495 1.085 8.495 1.415 8.435 1.415 8.435 1.085 8.085 1.085 8.085 1.415 8.025 1.415 8.025 1.085 7.675 1.085 7.675 1.415 7.615 1.415 7.615 1.085 7.265 1.085 7.265 1.415 7.205 1.415 7.205 1.085 6.855 1.085 6.855 1.415 6.795 1.415 6.795 1.085 6.445 1.085 6.445 1.415 6.385 1.415 6.385 1.085 6.08 1.085 6.08 1.11 6.035 1.11 6.035 1.415 5.975 1.415 5.975 1.05 6.02 1.05 6.02 0.66 5.885 0.66 5.885 0.475 5.945 0.475 5.945 0.6 6.14 0.6 6.14 0.73 6.08 0.73 6.08 1.025 6.385 1.025 6.385 0.615 6.295 0.615 6.295 0.475 6.355 0.475 6.355 0.555 6.705 0.555 6.705 0.475 6.765 0.475 6.765 0.615 6.445 0.615 6.445 1.025 7.205 1.025 7.205 0.615 7.115 0.615 7.115 0.475 7.175 0.475 7.175 0.555 7.525 0.555 7.525 0.475 7.585 0.475 7.585 0.615 7.265 0.615 7.265 1.025 8.345 1.025 8.345 0.615 7.935 0.615 7.935 0.475 7.995 0.475 7.995 0.555 8.345 0.555 8.345 0.475 8.405 0.475 8.405 1.025 9.62 1.025 9.62 0.615 8.755 0.615 8.755 0.475 8.815 0.475 8.815 0.555 9.165 0.555 9.165 0.475 9.225 0.475 9.225 0.555 9.575 0.555 9.575 0.475 9.68 0.475 9.68 1.025 9.725 1.025 ;
    END
  END Y
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0592 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2043 LAYER Metal1 ;
      ANTENNAMAXAREACAR 0.28977 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.68575625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.06 0.875 1.765 0.875 1.765 0.895 1.635 0.895 1.635 0.875 1.44 0.875 1.44 0.73 1.5 0.73 1.5 0.815 2 0.815 2 0.73 2.06 0.73 ;
    END
  END OE
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2916 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.436214 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.555 0.745 3.055 0.745 3.055 0.615 3.02 0.615 3.02 0.405 2.7 0.405 2.7 0.615 2.475 0.615 2.475 0.755 2.415 0.755 2.415 0.615 2.32 0.615 2.32 0.36 1.985 0.36 1.985 0.615 1.77 0.615 1.77 0.715 1.71 0.715 1.71 0.615 1.605 0.615 1.605 0.36 1.075 0.36 1.075 0.64 1 0.64 1 0.72 0.94 0.72 0.94 0.64 0.84 0.64 0.84 0.72 0.78 0.72 0.78 0.64 0.695 0.64 0.695 0.36 0.34 0.36 0.34 0.685 0.28 0.685 0.28 0.705 0.035 0.705 0.035 0.625 0.28 0.625 0.28 0.3 0.755 0.3 0.755 0.58 1.015 0.58 1.015 0.3 1.665 0.3 1.665 0.555 1.925 0.555 1.925 0.3 2.38 0.3 2.38 0.555 2.64 0.555 2.64 0.345 3.08 0.345 3.08 0.555 3.115 0.555 3.115 0.685 5.555 0.685 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 10 1.77 0 1.77 0 1.65 0.1 1.65 0.1 1.51 0.16 1.51 0.16 1.65 0.5 1.65 0.5 1.51 0.56 1.51 0.56 1.65 0.9 1.65 0.9 1.51 0.96 1.51 0.96 1.65 1.3 1.65 1.3 1.51 1.36 1.51 1.36 1.65 1.805 1.65 1.805 1.51 1.865 1.51 1.865 1.65 2.135 1.65 2.135 1.51 2.195 1.51 2.195 1.65 2.575 1.65 2.575 1.105 2.635 1.105 2.635 1.65 3.1 1.65 3.1 1.325 3.22 1.325 3.22 1.385 3.16 1.385 3.16 1.65 4 1.65 4 1.325 4.12 1.325 4.12 1.385 4.06 1.385 4.06 1.65 4.76 1.65 4.76 1.405 4.88 1.405 4.88 1.465 4.82 1.465 4.82 1.65 5.7 1.65 5.7 1.325 5.82 1.325 5.82 1.385 5.76 1.385 5.76 1.65 6.18 1.65 6.18 1.185 6.24 1.185 6.24 1.65 6.59 1.65 6.59 1.185 6.65 1.185 6.65 1.65 7 1.65 7 1.185 7.06 1.185 7.06 1.65 7.41 1.65 7.41 1.185 7.47 1.185 7.47 1.65 7.82 1.65 7.82 1.185 7.88 1.185 7.88 1.65 8.23 1.65 8.23 1.185 8.29 1.185 8.29 1.65 8.64 1.65 8.64 1.185 8.7 1.185 8.7 1.65 9.05 1.65 9.05 1.185 9.11 1.185 9.11 1.65 9.46 1.65 9.46 1.185 9.52 1.185 9.52 1.65 9.87 1.65 9.87 1.025 9.93 1.025 9.93 1.65 10 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 10 0.06 9.84 0.06 9.84 0.455 9.78 0.455 9.78 0.06 9.43 0.06 9.43 0.455 9.37 0.455 9.37 0.06 9.02 0.06 9.02 0.455 8.96 0.455 8.96 0.06 8.61 0.06 8.61 0.455 8.55 0.455 8.55 0.06 8.2 0.06 8.2 0.455 8.14 0.455 8.14 0.06 7.79 0.06 7.79 0.455 7.73 0.455 7.73 0.06 7.38 0.06 7.38 0.455 7.32 0.455 7.32 0.06 6.97 0.06 6.97 0.455 6.91 0.455 6.91 0.06 6.56 0.06 6.56 0.455 6.5 0.455 6.5 0.06 6.15 0.06 6.15 0.455 6.09 0.455 6.09 0.06 5.67 0.06 5.67 0.365 5.73 0.365 5.73 0.425 5.61 0.425 5.61 0.06 5.26 0.06 5.26 0.365 5.32 0.365 5.32 0.425 5.2 0.425 5.2 0.06 4.85 0.06 4.85 0.365 4.91 0.365 4.91 0.425 4.79 0.425 4.79 0.06 4.44 0.06 4.44 0.365 4.5 0.365 4.5 0.425 4.38 0.425 4.38 0.06 4.03 0.06 4.03 0.365 4.09 0.365 4.09 0.425 3.97 0.425 3.97 0.06 3.62 0.06 3.62 0.365 3.68 0.365 3.68 0.425 3.56 0.425 3.56 0.06 3.24 0.06 3.24 0.455 3.18 0.455 3.18 0.06 2.54 0.06 2.54 0.455 2.48 0.455 2.48 0.06 1.825 0.06 1.825 0.455 1.765 0.455 1.765 0.06 0.915 0.06 0.915 0.455 0.855 0.455 0.855 0.06 0.175 0.06 0.175 0.455 0.115 0.455 0.115 0.06 0 0.06 0 -0.06 10 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.92 0.95 5.875 0.95 5.875 1.225 5.6 1.225 5.6 1.305 4.25 1.305 4.25 1.225 2.735 1.225 2.735 1.005 2.43 1.005 2.43 1.225 2.37 1.225 2.37 1.035 2.03 1.035 2.03 1.12 1.97 1.12 1.97 1.06 1.63 1.06 1.63 1.12 1.57 1.12 1.57 1.06 1.125 1.06 1.125 1.12 1.065 1.12 1.065 1.06 0.725 1.06 0.725 1.12 0.665 1.12 0.665 1.06 0.325 1.06 0.325 1.225 0.265 1.225 0.265 0.9 0.325 0.9 0.325 1 0.44 1 0.44 0.46 0.56 0.46 0.56 0.52 0.5 0.52 0.5 1 1.28 1 1.28 0.46 1.4 0.46 1.4 0.52 1.34 0.52 1.34 1 1.865 1 1.865 0.975 2.16 0.975 2.16 0.52 2.085 0.52 2.085 0.46 2.22 0.46 2.22 0.975 2.37 0.975 2.37 0.945 2.795 0.945 2.795 1.165 4.31 1.165 4.31 1.245 5.54 1.245 5.54 1.165 5.815 1.165 5.815 0.89 5.86 0.89 5.86 0.83 5.92 0.83 ;
      POLYGON 5.76 0.765 5.715 0.765 5.715 1.065 5.29 1.065 5.29 1.145 5.23 1.145 5.23 1.065 4.47 1.065 4.47 1.145 4.41 1.145 4.41 1.065 3.66 1.065 3.66 1.005 5.655 1.005 5.655 0.585 3.385 0.585 3.385 0.43 3.445 0.43 3.445 0.525 3.795 0.525 3.795 0.43 3.855 0.43 3.855 0.525 4.205 0.525 4.205 0.43 4.265 0.43 4.265 0.525 4.615 0.525 4.615 0.43 4.675 0.43 4.675 0.525 5.025 0.525 5.025 0.43 5.085 0.43 5.085 0.525 5.435 0.525 5.435 0.43 5.495 0.43 5.495 0.525 5.715 0.525 5.715 0.645 5.76 0.645 ;
      POLYGON 5.18 0.905 2.955 0.905 2.955 1.02 2.895 1.02 2.895 0.775 2.8 0.775 2.8 0.505 2.92 0.505 2.92 0.715 2.955 0.715 2.955 0.845 5.18 0.845 ;
      POLYGON 1.18 0.9 0.6 0.9 0.6 0.74 0.68 0.74 0.68 0.82 1.1 0.82 1.1 0.74 1.18 0.74 ;
  END
END TBUFX20

MACRO TBUFX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX3 0 0 ;
  SIZE 2.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.2841 LAYER Metal1 ;
    ANTENNADIFFAREA 1.683175 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.117 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.97521375 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 84.79487175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.51 0.54 2.32 0.54 2.32 0.79 2.34 0.79 2.34 0.9 2.5 0.9 2.5 1.29 2.44 1.29 2.44 0.96 2.32 0.96 2.32 1.17 2.03 1.17 2.03 1.23 1.97 1.23 1.97 1.11 2.26 1.11 2.26 0.54 2.04 0.54 2.04 0.4 2.1 0.4 2.1 0.48 2.45 0.48 2.45 0.4 2.51 0.4 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 12.051282 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.735 0.69 1.675 0.69 1.675 0.33 0.895 0.33 0.895 0.815 0.965 0.815 0.965 0.895 0.835 0.895 0.835 0.89 0.44 0.89 0.44 0.83 0.835 0.83 0.835 0.27 1.735 0.27 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.25742575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.735 0.73 0.34 0.73 0.34 0.77 0.26 0.77 0.26 0.6 0.34 0.6 0.34 0.65 0.735 0.65 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 1.77 0 1.77 0 1.65 0.15 1.65 0.15 1.24 0.21 1.24 0.21 1.65 0.56 1.65 0.56 1.32 0.68 1.32 0.68 1.38 0.62 1.38 0.62 1.65 1.765 1.65 1.765 1.17 1.825 1.17 1.825 1.65 2.205 1.65 2.205 1.27 2.265 1.27 2.265 1.65 2.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.6 0.06 2.305 0.06 2.305 0.38 2.245 0.38 2.245 0.06 1.895 0.06 1.895 0.38 1.835 0.38 1.835 0.06 1.34 0.06 1.34 0.17 1.22 0.17 1.22 0.06 0.605 0.06 0.605 0.46 0.545 0.46 0.545 0.06 0 0.06 0 -0.06 2.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.105 1.01 1.66 1.01 1.66 1.22 0.415 1.22 0.415 1.36 0.355 1.36 0.355 1.05 0.1 1.05 0.1 0.44 0.205 0.44 0.205 0.38 0.265 0.38 0.265 0.5 0.16 0.5 0.16 0.99 0.415 0.99 0.415 1.16 1.6 1.16 1.6 0.95 2.045 0.95 2.045 0.705 2.105 0.705 ;
      POLYGON 1.94 0.85 1.5 0.85 1.5 1.02 1.44 1.02 1.44 0.79 1.445 0.79 1.445 0.43 1.575 0.43 1.575 0.49 1.505 0.49 1.505 0.79 1.88 0.79 1.88 0.56 1.94 0.56 ;
      POLYGON 1.345 0.65 1.125 0.65 1.125 1.06 0.795 1.06 0.795 1 1.065 1 1.065 0.57 0.995 0.57 0.995 0.51 1.125 0.51 1.125 0.59 1.345 0.59 ;
  END
END TBUFX3

MACRO TBUFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX4 0 0 ;
  SIZE 2.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3809 LAYER Metal1 ;
    ANTENNADIFFAREA 1.838675 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.14625 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.44205125 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 72.75897425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.515 1.33 2.455 1.33 2.455 1 2.12 1 2.12 1.15 2.105 1.15 2.105 1.33 2.045 1.33 2.045 1.09 2.06 1.09 2.06 0.55 1.945 0.55 1.945 0.41 2.005 0.41 2.005 0.49 2.355 0.49 2.355 0.41 2.415 0.41 2.415 0.55 2.12 0.55 2.12 0.79 2.14 0.79 2.14 0.94 2.515 0.94 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0585 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.6153845 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.64 0.67 1.52 0.67 1.52 0.61 1.58 0.61 1.58 0.34 0.895 0.34 0.895 0.625 0.965 0.625 0.965 0.705 0.895 0.705 0.895 0.89 0.445 0.89 0.445 0.83 0.835 0.83 0.835 0.28 1.64 0.28 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.2244225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.735 0.73 0.345 0.73 0.345 0.77 0.265 0.77 0.265 0.65 0.46 0.65 0.46 0.6 0.54 0.6 0.54 0.65 0.735 0.65 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 1.77 0 1.77 0 1.65 0.21 1.65 0.21 1.24 0.27 1.24 0.27 1.65 0.62 1.65 0.62 1.32 0.74 1.32 0.74 1.38 0.68 1.38 0.68 1.65 1.68 1.65 1.68 1.09 1.74 1.09 1.74 1.65 2.22 1.65 2.22 1.24 2.34 1.24 2.34 1.3 2.28 1.3 2.28 1.65 2.66 1.65 2.66 0.94 2.72 0.94 2.72 1.65 2.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.8 0.06 2.62 0.06 2.62 0.39 2.56 0.39 2.56 0.06 2.21 0.06 2.21 0.39 2.15 0.39 2.15 0.06 1.8 0.06 1.8 0.39 1.74 0.39 1.74 0.06 1.245 0.06 1.245 0.17 1.125 0.17 1.125 0.06 0.61 0.06 0.61 0.44 0.55 0.44 0.55 0.06 0 0.06 0 -0.06 2.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.96 0.99 1.58 0.99 1.58 1.22 0.475 1.22 0.475 1.36 0.415 1.36 0.415 1.05 0.105 1.05 0.105 0.49 0.21 0.49 0.21 0.43 0.27 0.43 0.27 0.55 0.165 0.55 0.165 0.99 0.475 0.99 0.475 1.16 1.52 1.16 1.52 0.93 1.9 0.93 1.9 0.745 1.96 0.745 ;
      POLYGON 1.8 0.83 1.42 0.83 1.42 1.06 1.36 1.06 1.36 0.44 1.48 0.44 1.48 0.5 1.42 0.5 1.42 0.77 1.74 0.77 1.74 0.595 1.8 0.595 ;
      POLYGON 1.26 0.785 1.125 0.785 1.125 1.06 0.86 1.06 0.86 1 1.065 1 1.065 0.525 0.995 0.525 0.995 0.465 1.125 0.465 1.125 0.725 1.26 0.725 ;
  END
END TBUFX4

MACRO TBUFX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX6 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4406 LAYER Metal1 ;
    ANTENNADIFFAREA 2.92225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.233775 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.439953 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 79.98716725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.18 0.59 4.13 0.59 4.13 1.29 4.07 1.29 4.07 0.96 3.72 0.96 3.72 1.29 3.66 1.29 3.66 0.96 3.52 0.96 3.52 1.05 3.31 1.05 3.31 1.29 3.25 1.29 3.25 0.99 3.46 0.99 3.46 0.64 3.3 0.64 3.3 0.45 3.36 0.45 3.36 0.58 3.52 0.58 3.52 0.79 3.54 0.79 3.54 0.9 4.07 0.9 4.07 0.59 3.71 0.59 3.71 0.45 3.77 0.45 3.77 0.53 4.12 0.53 4.12 0.45 4.18 0.45 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.11655 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.082368 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.03 0.325 2.89 0.325 2.89 0.33 1.39 0.33 1.39 0.92 0.59 0.92 0.59 0.86 0.635 0.86 0.635 0.815 0.765 0.815 0.765 0.86 1.33 0.86 1.33 0.27 2.83 0.27 2.83 0.265 3.03 0.265 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.074475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.5387715 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.23 0.76 1.17 0.76 1.17 0.715 0.985 0.715 0.985 0.755 0.865 0.755 0.865 0.715 0.34 0.715 0.34 0.92 0.22 0.92 0.22 0.86 0.26 0.86 0.26 0.655 1.17 0.655 1.17 0.64 1.23 0.64 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.77 0 1.77 0 1.65 0.12 1.65 0.12 1.18 0.18 1.18 0.18 1.65 0.545 1.65 0.545 1.18 0.605 1.18 0.605 1.65 0.955 1.65 0.955 1.18 1.015 1.18 1.015 1.65 1.365 1.65 1.365 1.54 1.485 1.54 1.485 1.65 2.2 1.65 2.2 1.2 2.32 1.2 2.32 1.26 2.26 1.26 2.26 1.65 3.045 1.65 3.045 1.03 3.105 1.03 3.105 1.65 3.455 1.65 3.455 1.17 3.515 1.17 3.515 1.65 3.865 1.65 3.865 1.06 3.925 1.06 3.925 1.65 4.275 1.65 4.275 0.9 4.335 0.9 4.335 1.65 4.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 0.06 4.385 0.06 4.385 0.43 4.325 0.43 4.325 0.06 3.975 0.06 3.975 0.43 3.915 0.43 3.915 0.06 3.565 0.06 3.565 0.43 3.505 0.43 3.505 0.06 3.19 0.06 3.19 0.485 3.065 0.485 3.065 0.425 3.13 0.425 3.13 0.06 2.73 0.06 2.73 0.17 2.61 0.17 2.61 0.06 2.235 0.06 2.235 0.17 2.115 0.17 2.115 0.06 1.74 0.06 1.74 0.17 1.62 0.17 1.62 0.06 1.19 0.06 1.19 0.54 1.13 0.54 1.13 0.06 0.49 0.06 0.49 0.335 0.55 0.335 0.55 0.395 0.43 0.395 0.43 0.06 0 0.06 0 -0.06 4.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.36 0.89 2.945 0.89 2.945 1.28 2.48 1.28 2.48 1.1 2.1 1.1 2.1 1.29 1.16 1.29 1.16 1.08 0.81 1.08 0.81 1.16 0.75 1.16 0.75 1.08 0.385 1.08 0.385 1.16 0.325 1.16 0.325 1.08 0.06 1.08 0.06 0.495 0.12 0.495 0.12 0.435 0.18 0.435 0.18 0.495 0.91 0.495 0.91 0.555 0.12 0.555 0.12 1.02 1.22 1.02 1.22 1.23 2.04 1.23 2.04 1.04 2.54 1.04 2.54 1.22 2.885 1.22 2.885 0.83 3.3 0.83 3.3 0.74 3.36 0.74 ;
      POLYGON 3.18 0.73 3.12 0.73 3.12 0.645 2.785 0.645 2.785 1.12 2.64 1.12 2.64 1.06 2.725 1.06 2.725 0.94 1.94 0.94 1.94 1.12 1.82 1.12 1.82 1.06 1.88 1.06 1.88 0.88 2.725 0.88 2.725 0.54 1.88 0.54 1.88 0.48 2.965 0.48 2.965 0.585 3.18 0.585 ;
      POLYGON 2.625 0.735 1.72 0.735 1.72 1.13 1.6 1.13 1.6 1.07 1.66 1.07 1.66 0.565 1.49 0.565 1.49 0.505 1.72 0.505 1.72 0.675 2.625 0.675 ;
  END
END TBUFX6

MACRO TBUFX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFX8 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.668 LAYER Metal1 ;
    ANTENNADIFFAREA 3.22625 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.292275 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.12838925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 70.1154735 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.59 0.59 4.54 0.59 4.54 1.29 4.48 1.29 4.48 0.96 4.13 0.96 4.13 1.29 4.07 1.29 4.07 0.96 3.72 0.96 3.72 1.29 3.66 1.29 3.66 0.96 3.52 0.96 3.52 1.05 3.31 1.05 3.31 1.29 3.25 1.29 3.25 0.99 3.46 0.99 3.46 0.64 3.3 0.64 3.3 0.45 3.36 0.45 3.36 0.58 3.52 0.58 3.52 0.79 3.54 0.79 3.54 0.9 4.48 0.9 4.48 0.59 3.71 0.59 3.71 0.45 3.77 0.45 3.77 0.53 4.12 0.53 4.12 0.45 4.18 0.45 4.18 0.53 4.53 0.53 4.53 0.45 4.59 0.45 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.11655 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.082368 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.03 0.325 2.89 0.325 2.89 0.33 1.39 0.33 1.39 0.92 0.59 0.92 0.59 0.86 0.635 0.86 0.635 0.815 0.765 0.815 0.765 0.86 1.33 0.86 1.33 0.27 2.83 0.27 2.83 0.265 3.03 0.265 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.074475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.5387715 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.23 0.76 1.17 0.76 1.17 0.715 0.985 0.715 0.985 0.755 0.865 0.755 0.865 0.715 0.34 0.715 0.34 0.92 0.22 0.92 0.22 0.86 0.26 0.86 0.26 0.655 1.17 0.655 1.17 0.64 1.23 0.64 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 1.77 0 1.77 0 1.65 0.12 1.65 0.12 1.18 0.18 1.18 0.18 1.65 0.545 1.65 0.545 1.18 0.605 1.18 0.605 1.65 0.955 1.65 0.955 1.18 1.015 1.18 1.015 1.65 1.365 1.65 1.365 1.54 1.485 1.54 1.485 1.65 2.2 1.65 2.2 1.2 2.32 1.2 2.32 1.26 2.26 1.26 2.26 1.65 3.045 1.65 3.045 1.03 3.105 1.03 3.105 1.65 3.455 1.65 3.455 1.17 3.515 1.17 3.515 1.65 3.865 1.65 3.865 1.06 3.925 1.06 3.925 1.65 4.275 1.65 4.275 1.06 4.335 1.06 4.335 1.65 4.685 1.65 4.685 0.9 4.745 0.9 4.745 1.65 5 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 0.06 4.795 0.06 4.795 0.43 4.735 0.43 4.735 0.06 4.385 0.06 4.385 0.43 4.325 0.43 4.325 0.06 3.975 0.06 3.975 0.43 3.915 0.43 3.915 0.06 3.565 0.06 3.565 0.43 3.505 0.43 3.505 0.06 3.19 0.06 3.19 0.485 3.065 0.485 3.065 0.425 3.13 0.425 3.13 0.06 2.73 0.06 2.73 0.17 2.61 0.17 2.61 0.06 2.235 0.06 2.235 0.17 2.115 0.17 2.115 0.06 1.74 0.06 1.74 0.17 1.62 0.17 1.62 0.06 1.19 0.06 1.19 0.54 1.13 0.54 1.13 0.06 0.49 0.06 0.49 0.335 0.55 0.335 0.55 0.395 0.43 0.395 0.43 0.06 0 0.06 0 -0.06 5 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.36 0.89 2.945 0.89 2.945 1.28 2.48 1.28 2.48 1.1 2.1 1.1 2.1 1.29 1.16 1.29 1.16 1.08 0.81 1.08 0.81 1.16 0.75 1.16 0.75 1.08 0.385 1.08 0.385 1.16 0.325 1.16 0.325 1.08 0.06 1.08 0.06 0.495 0.12 0.495 0.12 0.435 0.18 0.435 0.18 0.495 0.91 0.495 0.91 0.555 0.12 0.555 0.12 1.02 1.22 1.02 1.22 1.23 2.04 1.23 2.04 1.04 2.54 1.04 2.54 1.22 2.885 1.22 2.885 0.83 3.3 0.83 3.3 0.74 3.36 0.74 ;
      POLYGON 3.18 0.73 3.12 0.73 3.12 0.645 2.785 0.645 2.785 1.12 2.64 1.12 2.64 1.06 2.725 1.06 2.725 0.94 1.94 0.94 1.94 1.12 1.82 1.12 1.82 1.06 1.88 1.06 1.88 0.88 2.725 0.88 2.725 0.54 1.88 0.54 1.88 0.48 2.965 0.48 2.965 0.585 3.18 0.585 ;
      POLYGON 2.625 0.735 1.66 0.735 1.66 1.07 1.72 1.07 1.72 1.13 1.6 1.13 1.6 0.565 1.49 0.565 1.49 0.505 1.66 0.505 1.66 0.675 2.625 0.675 ;
  END
END TBUFX8

MACRO TBUFXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TBUFXL 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.9075 LAYER Metal1 ;
    ANTENNADIFFAREA 1.080725 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXAREACAR 28.00925925 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 216.388889 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.745 1.11 1.66 1.11 1.66 0.98 1.685 0.98 1.685 0.605 1.675 0.605 1.675 0.485 1.735 0.485 1.735 0.565 1.745 0.565 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 19.72222225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.415 0.365 0.685 0.365 0.685 0.625 0.845 0.625 0.845 1.025 0.565 1.025 0.565 1.085 0.435 1.085 0.435 1.025 0.385 1.025 0.385 0.965 0.785 0.965 0.785 0.685 0.625 0.685 0.625 0.305 1.415 0.305 ;
    END
  END A
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.9444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.685 0.865 0.2 0.865 0.2 0.745 0.26 0.745 0.26 0.6 0.34 0.6 0.34 0.785 0.685 0.785 ;
    END
  END OE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.285 0.13 1.285 0.13 1.65 0.48 1.65 0.48 1.54 0.6 1.54 0.6 1.65 1.45 1.65 1.45 1.51 1.51 1.51 1.51 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.575 0.06 1.575 0.52 1.53 0.52 1.53 0.58 1.47 0.58 1.47 0.46 1.515 0.46 1.515 0.06 1.105 0.06 1.105 0.17 0.985 0.17 0.985 0.06 0.525 0.06 0.525 0.5 0.465 0.5 0.465 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.67 1.435 1.61 1.435 1.61 1.375 1.35 1.375 1.35 1.44 0.275 1.44 0.275 1.185 0.04 1.185 0.04 0.52 0.1 0.52 0.1 0.46 0.16 0.46 0.16 0.58 0.1 0.58 0.1 1.125 0.335 1.125 0.335 1.38 1.29 1.38 1.29 1.315 1.67 1.315 ;
      POLYGON 1.585 0.74 1.36 0.74 1.36 0.895 1.17 0.895 1.17 1.06 1.11 1.06 1.11 0.835 1.3 0.835 1.3 0.575 1.22 0.575 1.22 0.515 1.36 0.515 1.36 0.68 1.585 0.68 ;
      POLYGON 1.2 0.735 1.005 0.735 1.005 1.28 0.715 1.28 0.715 1.22 0.945 1.22 0.945 0.525 0.785 0.525 0.785 0.465 1.005 0.465 1.005 0.675 1.2 0.675 ;
  END
END TBUFXL

MACRO TIEHI
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIEHI 0 0 ;
  SIZE 0.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.117 LAYER Metal1 ;
    ANTENNADIFFAREA 0.1812 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.9 0.14 1.4 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 1.77 0 1.77 0 1.65 0.275 1.65 0.275 0.9 0.335 0.9 0.335 1.65 0.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 0.06 0.335 0.06 0.335 0.49 0.275 0.49 0.275 0.06 0 0.06 0 -0.06 0.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.205 0.8 0.125 0.8 0.125 0.65 0.07 0.65 0.07 0.355 0.15 0.355 0.15 0.57 0.205 0.57 ;
  END
END TIEHI

MACRO TIELO
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIELO 0 0 ;
  SIZE 0.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0996 LAYER Metal1 ;
    ANTENNADIFFAREA 0.1448 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.16 0.14 0.66 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 1.77 0 1.77 0 1.65 0.275 1.65 0.275 0.95 0.335 0.95 0.335 1.65 0.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.6 0.06 0.335 0.06 0.335 0.52 0.275 0.52 0.275 0.06 0 0.06 0 -0.06 0.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 0.225 0.85 0.15 0.85 0.15 1.29 0.07 1.29 0.07 0.77 0.225 0.77 ;
  END
END TIELO

MACRO TLATNCAX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX12 0 0 ;
  SIZE 5.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.1963 LAYER Metal1 ;
    ANTENNADIFFAREA 4.086825 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.62055 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.15075325 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 40.826686 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.34 0.99 0.67 0.99 0.67 1.02 0.61 1.02 0.61 0.9 0.99 0.9 0.99 0.57 0.61 0.57 0.61 0.26 0.67 0.26 0.67 0.51 1.02 0.51 1.02 0.26 1.08 0.26 1.08 0.51 1.43 0.51 1.43 0.26 1.49 0.26 1.49 0.51 1.84 0.51 1.84 0.26 1.9 0.26 1.9 0.51 2.25 0.51 2.25 0.26 2.31 0.26 2.31 0.57 1.05 0.57 1.05 0.79 1.14 0.79 1.14 0.93 2.34 0.93 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.34 1.22 5.26 1.22 5.26 1.06 5.13 1.06 5.13 0.85 5.21 0.85 5.21 0.98 5.34 0.98 ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.51 0.895 0.235 0.895 0.235 0.7 0.205 0.7 0.205 0.62 0.325 0.62 0.325 0.815 0.51 0.815 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 1.77 0 1.77 0 1.65 0.375 1.65 0.375 1.285 0.435 1.285 0.435 1.65 0.785 1.65 0.785 1.28 0.905 1.28 0.905 1.34 0.845 1.34 0.845 1.65 1.195 1.65 1.195 1.28 1.315 1.28 1.315 1.34 1.255 1.34 1.255 1.65 1.605 1.65 1.605 1.28 1.725 1.28 1.725 1.34 1.665 1.34 1.665 1.65 2.015 1.65 2.015 1.28 2.135 1.28 2.135 1.34 2.075 1.34 2.075 1.65 2.455 1.65 2.455 1.41 2.575 1.41 2.575 1.47 2.515 1.47 2.515 1.65 2.84 1.65 2.84 1.41 2.96 1.41 2.96 1.47 2.9 1.47 2.9 1.65 3.31 1.65 3.31 1.41 3.43 1.41 3.43 1.47 3.37 1.47 3.37 1.65 3.78 1.65 3.78 1.41 3.9 1.41 3.9 1.47 3.84 1.47 3.84 1.65 4.28 1.65 4.28 1.51 4.34 1.51 4.34 1.65 5.235 1.65 5.235 1.32 5.295 1.32 5.295 1.65 5.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.6 0.06 5.325 0.06 5.325 0.43 5.205 0.43 5.205 0.37 5.265 0.37 5.265 0.06 4.285 0.06 4.285 0.52 4.225 0.52 4.225 0.06 3.34 0.06 3.34 0.43 3.4 0.43 3.4 0.49 3.28 0.49 3.28 0.06 2.515 0.06 2.515 0.57 2.455 0.57 2.455 0.06 2.105 0.06 2.105 0.38 2.045 0.38 2.045 0.06 1.695 0.06 1.695 0.38 1.635 0.38 1.635 0.06 1.285 0.06 1.285 0.38 1.225 0.38 1.225 0.06 0.875 0.06 0.875 0.38 0.815 0.38 0.815 0.06 0.465 0.06 0.465 0.52 0.405 0.52 0.405 0.06 0 0.06 0 -0.06 5.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.53 1.44 5.47 1.44 5.47 0.59 5.045 0.59 5.045 0.41 4.445 0.41 4.445 0.81 4.275 0.81 4.275 0.815 4.155 0.815 4.155 0.81 3.415 0.81 3.415 0.75 4.385 0.75 4.385 0.35 5.105 0.35 5.105 0.53 5.44 0.53 5.44 0.47 5.53 0.47 ;
      POLYGON 5.37 0.81 5.31 0.81 5.31 0.75 5.03 0.75 5.03 1.14 4.79 1.14 4.79 1.08 4.97 1.08 4.97 0.75 4.885 0.75 4.885 0.57 4.59 0.57 4.59 0.51 4.945 0.51 4.945 0.69 5.37 0.69 ;
      POLYGON 4.87 0.975 2.835 0.975 2.835 0.99 2.66 0.99 2.66 0.93 2.775 0.93 2.775 0.45 2.835 0.45 2.835 0.915 3.675 0.915 3.675 0.91 3.795 0.91 3.795 0.915 4.545 0.915 4.545 0.83 4.605 0.83 4.605 0.915 4.81 0.915 4.81 0.855 4.87 0.855 ;
      POLYGON 4.7 1.425 4.63 1.425 4.63 1.31 2.235 1.31 2.235 1.18 0.075 1.18 0.075 0.86 0.045 0.86 0.045 0.485 0.07 0.485 0.07 0.425 0.13 0.425 0.13 0.545 0.105 0.545 0.105 0.8 0.135 0.8 0.135 1.12 2.295 1.12 2.295 1.25 4.69 1.25 4.69 1.305 4.7 1.305 ;
      POLYGON 4.135 1.15 2.5 1.15 2.5 0.73 2.155 0.73 2.155 0.67 2.615 0.67 2.615 0.29 2.995 0.29 2.995 0.43 3.09 0.43 3.09 0.59 3.5 0.59 3.5 0.57 3.77 0.57 3.77 0.63 3.55 0.63 3.55 0.65 3.03 0.65 3.03 0.49 2.935 0.49 2.935 0.35 2.675 0.35 2.675 0.73 2.56 0.73 2.56 1.09 4.135 1.09 ;
  END
END TLATNCAX12

MACRO TLATNCAX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX16 0 0 ;
  SIZE 7.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.998175 LAYER Metal1 ;
    ANTENNADIFFAREA 5.280575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.81135 LAYER Metal1 ;
      ANTENNAMAXAREACAR 4.9278055 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 38.90552775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.215 0.63 3.125 0.63 3.125 0.645 2.775 0.645 2.775 1.01 3.16 1.01 3.16 1.07 0.58 1.07 0.58 1.01 0.665 1.01 0.665 0.54 0.725 0.54 0.725 1.01 1.045 1.01 1.045 0.57 1.165 0.57 1.165 0.63 1.105 0.63 1.105 1.01 1.455 1.01 1.455 0.57 1.575 0.57 1.575 0.63 1.515 0.63 1.515 1.01 1.865 1.01 1.865 0.57 1.985 0.57 1.985 0.63 1.93 0.63 1.93 1.01 2.26 1.01 2.26 0.57 2.395 0.57 2.395 0.63 2.32 0.63 2.32 0.79 2.34 0.79 2.34 1.01 2.715 1.01 2.715 0.525 2.775 0.525 2.775 0.585 3.08 0.585 3.08 0.57 3.215 0.57 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.5185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 6.66 0.67 6.78 1.01 ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 0.73 0.41 0.73 0.41 0.97 0.33 0.97 0.33 0.65 0.46 0.65 0.46 0.6 0.54 0.6 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 1.77 0 1.77 0 1.65 0.375 1.65 0.375 1.335 0.495 1.335 0.495 1.395 0.435 1.395 0.435 1.65 0.785 1.65 0.785 1.335 0.905 1.335 0.905 1.395 0.845 1.395 0.845 1.65 1.195 1.65 1.195 1.335 1.315 1.335 1.315 1.395 1.255 1.395 1.255 1.65 1.605 1.65 1.605 1.335 1.725 1.335 1.725 1.395 1.665 1.395 1.665 1.65 2.015 1.65 2.015 1.335 2.135 1.335 2.135 1.395 2.075 1.395 2.075 1.65 2.425 1.65 2.425 1.335 2.545 1.335 2.545 1.395 2.485 1.395 2.485 1.65 2.835 1.65 2.835 1.335 2.955 1.335 2.955 1.395 2.895 1.395 2.895 1.65 3.245 1.65 3.245 1.335 3.365 1.335 3.365 1.395 3.305 1.395 3.305 1.65 3.72 1.65 3.72 1.335 3.84 1.335 3.84 1.395 3.78 1.395 3.78 1.65 4.19 1.65 4.19 1.335 4.31 1.335 4.31 1.395 4.25 1.395 4.25 1.65 4.66 1.65 4.66 1.335 4.78 1.335 4.78 1.395 4.72 1.395 4.72 1.65 5.16 1.65 5.16 1.51 5.22 1.51 5.22 1.65 5.555 1.65 5.555 1.365 5.675 1.365 5.675 1.425 5.615 1.425 5.615 1.65 6.765 1.65 6.765 1.11 6.825 1.11 6.825 1.65 7.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.2 0.06 6.885 0.06 6.885 0.25 6.765 0.25 6.765 0.19 6.825 0.19 6.825 0.06 5.73 0.06 5.73 0.2 5.67 0.2 5.67 0.06 5.09 0.06 5.09 0.485 5.03 0.485 5.03 0.06 4.25 0.06 4.25 0.315 4.31 0.315 4.31 0.375 4.19 0.375 4.19 0.06 3.415 0.06 3.415 0.485 3.355 0.485 3.355 0.06 2.98 0.06 2.98 0.485 2.92 0.485 2.92 0.06 2.57 0.06 2.57 0.485 2.51 0.485 2.51 0.06 2.16 0.06 2.16 0.485 2.1 0.485 2.1 0.06 1.75 0.06 1.75 0.485 1.69 0.485 1.69 0.06 1.34 0.06 1.34 0.485 1.28 0.485 1.28 0.06 0.93 0.06 0.93 0.485 0.87 0.485 0.87 0.06 0.52 0.06 0.52 0.485 0.46 0.485 0.46 0.06 0 0.06 0 -0.06 7.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.1 0.96 7.07 0.96 7.07 1.135 7.01 1.135 7.01 0.9 7.04 0.9 7.04 0.41 6.605 0.41 6.605 0.405 5.25 0.405 5.25 0.695 4.61 0.695 4.61 0.755 4.49 0.755 4.49 0.695 4.01 0.695 4.01 0.755 3.89 0.755 3.89 0.635 5.19 0.635 5.19 0.345 6.665 0.345 6.665 0.35 7.1 0.35 ;
      POLYGON 6.94 0.82 6.88 0.82 6.88 0.57 6.54 0.57 6.54 1.265 4.88 1.265 4.88 1.235 0.17 1.235 0.17 0.54 0.23 0.54 0.23 1.175 4.94 1.175 4.94 1.205 6.48 1.205 6.48 0.94 6.085 0.94 6.085 0.82 6.145 0.82 6.145 0.88 6.48 0.88 6.48 0.51 6.94 0.51 ;
      POLYGON 6.38 0.625 5.985 0.625 5.985 1.045 6.165 1.045 6.165 1.105 5.925 1.105 5.925 0.945 5.51 0.945 5.51 0.81 5.57 0.81 5.57 0.885 5.925 0.885 5.925 0.565 6.32 0.565 6.32 0.505 6.38 0.505 ;
      POLYGON 5.825 0.785 5.765 0.785 5.765 0.71 5.41 0.71 5.41 1.1 5.35 1.1 5.35 0.915 3.475 0.915 3.475 0.795 3.535 0.795 3.535 0.855 4.115 0.855 4.115 0.795 4.175 0.795 4.175 0.855 4.99 0.855 4.99 0.795 5.05 0.795 5.05 0.855 5.35 0.855 5.35 0.505 5.41 0.505 5.41 0.65 5.825 0.65 ;
      POLYGON 5.015 1.075 3.315 1.075 3.315 0.815 3.08 0.815 3.08 0.755 3.315 0.755 3.315 0.635 3.72 0.635 3.72 0.475 4.75 0.475 4.75 0.535 3.78 0.535 3.78 0.695 3.375 0.695 3.375 1.015 5.015 1.015 ;
  END
END TLATNCAX16

MACRO TLATNCAX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX2 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.5861 LAYER Metal1 ;
    ANTENNADIFFAREA 1.92825 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1719 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.226876 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 71.69284475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.75 1.02 0.67 1.02 0.67 0.73 0.66 0.73 0.66 0.52 0.74 0.52 0.74 0.68 0.75 0.68 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.81 0.935 2.695 0.935 2.695 1.055 2.615 1.055 2.615 0.67 2.695 0.67 2.695 0.815 2.81 0.815 ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 0.73 0.46 0.73 0.46 1.02 0.38 1.02 0.38 0.65 0.46 0.65 0.46 0.6 0.54 0.6 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 1.77 0 1.77 0 1.65 0.455 1.65 0.455 1.28 0.515 1.28 0.515 1.65 0.895 1.65 0.895 1.41 1.015 1.41 1.015 1.47 0.955 1.47 0.955 1.65 1.355 1.65 1.355 1.51 1.415 1.51 1.415 1.65 1.825 1.65 1.825 1.51 1.885 1.51 1.885 1.65 2.68 1.65 2.68 1.155 2.74 1.155 2.74 1.65 3.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 0.06 2.74 0.06 2.74 0.19 2.8 0.19 2.8 0.25 2.68 0.25 2.68 0.06 1.785 0.06 1.785 0.2 1.725 0.2 1.725 0.06 0.925 0.06 0.925 0.5 0.865 0.5 0.865 0.06 0.515 0.06 0.515 0.5 0.455 0.5 0.455 0.06 0 0.06 0 -0.06 3.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.13 1.15 2.955 1.15 2.955 1.09 3.07 1.09 3.07 0.41 1.885 0.41 1.885 0.35 3.13 0.35 ;
      POLYGON 2.97 0.825 2.91 0.825 2.91 0.57 2.515 0.57 2.515 1.15 2.275 1.15 2.275 1.09 2.455 1.09 2.455 0.63 2.19 0.63 2.19 0.51 2.97 0.51 ;
      POLYGON 2.355 0.985 2.295 0.985 2.295 0.925 1.305 0.925 1.305 0.99 1.185 0.99 1.185 0.52 1.245 0.52 1.245 0.865 2.03 0.865 2.03 0.76 2.09 0.76 2.09 0.865 2.355 0.865 ;
      POLYGON 2.185 1.435 2.125 1.435 2.125 1.31 0.615 1.31 0.615 1.18 0.22 1.18 0.22 0.52 0.28 0.52 0.28 1.12 0.675 1.12 0.675 1.25 2.185 1.25 ;
      POLYGON 1.68 1.15 1.025 1.15 1.025 0.83 0.85 0.83 0.85 0.77 1.025 0.77 1.025 0.36 1.445 0.36 1.445 0.63 1.385 0.63 1.385 0.42 1.085 0.42 1.085 1.09 1.68 1.09 ;
  END
END TLATNCAX2

MACRO TLATNCAX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX20 0 0 ;
  SIZE 8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.79815 LAYER Metal1 ;
    ANTENNADIFFAREA 5.94835 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0008 LAYER Metal1 ;
      ANTENNAMAXAREACAR 4.7943145 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 38.49220625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.83 1.4 7.77 1.4 7.77 0.845 7.42 0.845 7.42 1.405 7.36 1.405 7.36 0.845 7.01 0.845 7.01 1.405 6.95 1.405 6.95 0.845 6.6 0.845 6.6 1.405 6.54 1.405 6.54 0.845 6.19 0.845 6.19 1.405 6.13 1.405 6.13 0.845 5.78 0.845 5.78 1.405 5.72 1.405 5.72 0.845 5.37 0.845 5.37 1.405 5.31 1.405 5.31 0.845 4.96 0.845 4.96 1.405 4.9 1.405 4.9 0.845 4.55 0.845 4.55 1.405 4.49 1.405 4.49 0.92 4.46 0.92 4.46 0.355 4.52 0.355 4.52 0.785 4.87 0.785 4.87 0.355 4.93 0.355 4.93 0.785 5.235 0.785 5.235 0.6 5.28 0.6 5.28 0.355 5.34 0.355 5.34 0.66 5.295 0.66 5.295 0.785 5.69 0.785 5.69 0.355 5.75 0.355 5.75 0.785 6.055 0.785 6.055 0.625 6.1 0.625 6.1 0.355 6.16 0.355 6.16 0.685 6.115 0.685 6.115 0.785 6.51 0.785 6.51 0.355 6.57 0.355 6.57 0.785 6.875 0.785 6.875 0.6 6.92 0.6 6.92 0.355 6.98 0.355 6.98 0.66 6.935 0.66 6.935 0.785 7.33 0.785 7.33 0.355 7.39 0.355 7.39 0.785 7.695 0.785 7.695 0.6 7.74 0.6 7.74 0.355 7.8 0.355 7.8 0.66 7.755 0.66 7.755 0.785 7.83 0.785 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.61 0.54 1.11 ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.61 0.34 1.11 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 1.77 0 1.77 0 1.65 0.405 1.65 0.405 1.21 0.465 1.21 0.465 1.65 1.18 1.65 1.18 1.41 1.3 1.41 1.3 1.47 1.24 1.47 1.24 1.65 1.65 1.65 1.65 1.49 1.77 1.49 1.77 1.55 1.71 1.55 1.71 1.65 2.09 1.65 2.09 1.285 2.15 1.285 2.15 1.65 2.5 1.65 2.5 1.185 2.56 1.185 2.56 1.65 2.91 1.65 2.91 1.185 2.97 1.185 2.97 1.65 3.32 1.65 3.32 1.185 3.38 1.185 3.38 1.65 3.875 1.65 3.875 1.185 3.935 1.185 3.935 1.65 4.285 1.65 4.285 1.185 4.345 1.185 4.345 1.65 4.695 1.65 4.695 0.945 4.755 0.945 4.755 1.65 5.105 1.65 5.105 0.945 5.165 0.945 5.165 1.65 5.515 1.65 5.515 0.945 5.575 0.945 5.575 1.65 5.925 1.65 5.925 0.945 5.985 0.945 5.985 1.65 6.335 1.65 6.335 0.945 6.395 0.945 6.395 1.65 6.745 1.65 6.745 0.945 6.805 0.945 6.805 1.65 7.155 1.65 7.155 0.945 7.215 0.945 7.215 1.65 7.565 1.65 7.565 0.945 7.625 0.945 7.625 1.65 8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8 0.06 7.595 0.06 7.595 0.66 7.535 0.66 7.535 0.06 7.185 0.06 7.185 0.66 7.125 0.66 7.125 0.06 6.775 0.06 6.775 0.66 6.715 0.66 6.715 0.06 6.365 0.06 6.365 0.66 6.305 0.66 6.305 0.06 5.955 0.06 5.955 0.66 5.895 0.66 5.895 0.06 5.545 0.06 5.545 0.66 5.485 0.66 5.485 0.06 5.135 0.06 5.135 0.66 5.075 0.66 5.075 0.06 4.725 0.06 4.725 0.66 4.665 0.66 4.665 0.06 4.295 0.06 4.295 0.475 4.235 0.475 4.235 0.06 3.35 0.06 3.35 0.385 3.41 0.385 3.41 0.445 3.29 0.445 3.29 0.06 2.63 0.06 2.63 0.385 2.69 0.385 2.69 0.445 2.57 0.445 2.57 0.06 1.8 0.06 1.8 0.17 1.68 0.17 1.68 0.06 1.33 0.06 1.33 0.17 1.21 0.17 1.21 0.06 0.455 0.06 0.455 0.35 0.395 0.35 0.395 0.06 0 0.06 0 -0.06 8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.36 1.085 4.14 1.085 4.14 1.405 4.08 1.405 4.08 1.085 3.73 1.085 3.73 1.405 3.67 1.405 3.67 1.085 3.175 1.085 3.175 1.405 3.115 1.405 3.115 1.085 2.765 1.085 2.765 1.405 2.705 1.405 2.705 1.085 2.355 1.085 2.355 1.405 2.295 1.405 2.295 1.025 4.3 1.025 4.3 0.76 4.075 0.76 4.075 0.605 2.33 0.605 2.33 0.585 2.26 0.585 2.26 0.525 2.38 0.525 2.38 0.545 2.88 0.545 2.88 0.525 3 0.525 3 0.545 3.875 0.545 3.875 0.485 3.935 0.485 3.935 0.545 4.135 0.545 4.135 0.7 4.36 0.7 ;
      POLYGON 4.2 0.925 2.165 0.925 2.165 1.15 1.725 1.15 1.725 1.04 1.445 1.04 1.445 0.92 1.505 0.92 1.505 0.63 1.12 0.63 1.12 0.57 1.565 0.57 1.565 0.98 1.785 0.98 1.785 1.09 2.105 1.09 2.105 0.865 4.2 0.865 ;
      POLYGON 3.835 0.765 2.005 0.765 2.005 0.99 1.885 0.99 1.885 0.93 1.945 0.93 1.945 0.47 1.02 0.47 1.02 0.545 0.96 0.545 0.96 0.41 2.005 0.41 2.005 0.705 3.835 0.705 ;
      POLYGON 1.93 1.31 1.08 1.31 1.08 1.395 0.995 1.395 0.995 1.5 0.935 1.5 0.935 1.395 0.64 1.395 0.64 0.51 0.16 0.51 0.16 1.21 0.26 1.21 0.26 1.33 0.2 1.33 0.2 1.27 0.1 1.27 0.1 0.45 0.19 0.45 0.19 0.255 0.25 0.255 0.25 0.45 0.7 0.45 0.7 1.335 1.02 1.335 1.02 1.25 1.93 1.25 ;
      POLYGON 1.405 0.82 0.92 0.82 0.92 1.235 0.86 1.235 0.86 0.85 0.8 0.85 0.8 0.255 0.86 0.255 0.86 0.76 1.405 0.76 ;
  END
END TLATNCAX20

MACRO TLATNCAX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX3 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8082 LAYER Metal1 ;
    ANTENNADIFFAREA 1.982975 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.22725 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.95687575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 62.87788775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.31 0.68 2.92 0.68 2.92 0.79 2.94 0.79 2.94 1.01 3.31 1.01 3.31 1.4 3.25 1.4 3.25 1.07 2.9 1.07 2.9 1.4 2.84 1.4 2.84 1.01 2.86 1.01 2.86 0.66 2.84 0.66 2.84 0.54 2.92 0.54 2.92 0.62 3.25 0.62 3.25 0.54 3.31 0.54 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.855 1.03 0.775 1.03 0.775 0.895 0.49 0.895 0.49 0.815 0.855 0.815 ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.23 0.82 0.15 0.82 0.15 0.54 0.06 0.54 0.06 0.41 0.14 0.41 0.14 0.46 0.23 0.46 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 1.77 0 1.77 0 1.65 0.125 1.65 0.125 0.995 0.185 0.995 0.185 1.65 0.765 1.65 0.765 1.29 0.825 1.29 0.825 1.65 1.57 1.65 1.57 1.29 1.63 1.29 1.63 1.65 2.195 1.65 2.195 1.31 2.315 1.31 2.315 1.37 2.255 1.37 2.255 1.65 2.635 1.65 2.635 1.28 2.695 1.28 2.695 1.65 3.045 1.65 3.045 1.17 3.105 1.17 3.105 1.65 3.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 0.06 3.105 0.06 3.105 0.52 3.045 0.52 3.045 0.06 2.665 0.06 2.665 0.43 2.725 0.43 2.725 0.49 2.605 0.49 2.605 0.06 1.715 0.06 1.715 0.2 1.655 0.2 1.655 0.06 0.91 0.06 0.91 0.395 0.85 0.395 0.85 0.06 0.225 0.06 0.225 0.2 0.165 0.2 0.165 0.06 0 0.06 0 -0.06 3.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.74 0.82 2.725 0.82 2.725 1.135 2.49 1.135 2.49 1.4 2.43 1.4 2.43 1.075 2.665 1.075 2.665 0.65 2.365 0.65 2.365 0.63 2.295 0.63 2.295 0.57 2.415 0.57 2.415 0.59 2.725 0.59 2.725 0.7 2.74 0.7 ;
      POLYGON 2.565 0.975 1.835 0.975 1.835 1.315 1.775 1.315 1.775 0.975 1.465 0.975 1.465 0.915 1.975 0.915 1.975 0.455 2.035 0.455 2.035 0.915 2.505 0.915 2.505 0.84 2.565 0.84 ;
      POLYGON 2.38 0.815 2.235 0.815 2.235 0.79 2.135 0.79 2.135 0.355 1.875 0.355 1.875 0.36 1.505 0.36 1.505 0.32 1.185 0.32 1.185 1.025 1.015 1.025 1.015 1.19 0.62 1.19 0.62 1.315 0.56 1.315 0.56 1.13 0.955 1.13 0.955 0.965 1.125 0.965 1.125 0.555 0.665 0.555 0.665 0.545 0.585 0.545 0.585 0.485 0.705 0.485 0.705 0.495 1.125 0.495 1.125 0.26 1.36 0.26 1.36 0.24 1.48 0.24 1.48 0.26 1.565 0.26 1.565 0.3 1.815 0.3 1.815 0.295 2.195 0.295 2.195 0.73 2.295 0.73 2.295 0.755 2.38 0.755 ;
      POLYGON 1.84 0.73 1.345 0.73 1.345 1.255 1.175 1.255 1.175 1.315 1.115 1.315 1.115 1.195 1.285 1.195 1.285 0.485 1.405 0.485 1.405 0.545 1.345 0.545 1.345 0.67 1.84 0.67 ;
      POLYGON 1.025 0.865 0.965 0.865 0.965 0.715 0.39 0.715 0.39 1.02 0.33 1.02 0.33 0.54 0.39 0.54 0.39 0.655 1.025 0.655 ;
  END
END TLATNCAX3

MACRO TLATNCAX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX4 0 0 ;
  SIZE 3.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8063 LAYER Metal1 ;
    ANTENNADIFFAREA 2.243375 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2565 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.04210525 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 56.6842105 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.2 0.99 1.08 0.99 1.08 0.96 0.7 0.96 0.7 1.02 0.64 1.02 0.64 0.9 0.66 0.9 0.66 0.51 0.72 0.51 0.72 0.57 1.055 0.57 1.055 0.55 1.175 0.55 1.175 0.61 1.105 0.61 1.105 0.63 0.72 0.63 0.72 0.79 0.74 0.79 0.74 0.9 1.14 0.9 1.14 0.93 1.2 0.93 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.25 0.895 3.03 0.895 3.03 1.06 2.95 1.06 2.95 0.78 3.25 0.78 ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 0.73 0.41 0.73 0.41 0.97 0.33 0.97 0.33 0.65 0.46 0.65 0.46 0.6 0.54 0.6 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 1.77 0 1.77 0 1.65 0.405 1.65 0.405 1.28 0.465 1.28 0.465 1.65 0.845 1.65 0.845 1.28 0.965 1.28 0.965 1.34 0.905 1.34 0.905 1.65 1.345 1.65 1.345 1.51 1.405 1.51 1.405 1.65 1.78 1.65 1.78 1.51 1.84 1.51 1.84 1.65 2.22 1.65 2.22 1.41 2.34 1.41 2.34 1.47 2.28 1.47 2.28 1.65 3.015 1.65 3.015 1.16 3.075 1.16 3.075 1.65 3.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 0.06 3.135 0.06 3.135 0.36 3.015 0.36 3.015 0.3 3.075 0.3 3.075 0.06 2.12 0.06 2.12 0.425 2.18 0.425 2.18 0.545 2.12 0.545 2.12 0.485 2.06 0.485 2.06 0.06 1.35 0.06 1.35 0.5 1.29 0.5 1.29 0.06 0.895 0.06 0.895 0.41 0.955 0.41 0.955 0.47 0.835 0.47 0.835 0.06 0.515 0.06 0.515 0.5 0.455 0.5 0.455 0.06 0 0.06 0 -0.06 3.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.57 1.155 3.25 1.155 3.25 1.095 3.51 1.095 3.51 0.52 2.855 0.52 2.855 0.325 2.22 0.325 2.22 0.265 2.915 0.265 2.915 0.46 3.28 0.46 3.28 0.4 3.34 0.4 3.34 0.46 3.57 0.46 ;
      POLYGON 3.41 0.74 3.35 0.74 3.35 0.68 2.85 0.68 2.85 1.155 2.6 1.155 2.6 1.095 2.79 1.095 2.79 0.68 2.525 0.68 2.525 0.425 2.585 0.425 2.585 0.62 3.41 0.62 ;
      POLYGON 2.69 0.98 2.63 0.98 2.63 0.88 1.73 0.88 1.73 0.99 1.61 0.99 1.61 0.93 1.67 0.93 1.67 0.83 1.61 0.83 1.61 0.52 1.67 0.52 1.67 0.77 1.73 0.77 1.73 0.82 2.365 0.82 2.365 0.76 2.425 0.76 2.425 0.82 2.69 0.82 ;
      POLYGON 2.595 1.44 2.535 1.44 2.535 1.315 2.44 1.315 2.44 1.31 1.065 1.31 1.065 1.18 0.17 1.18 0.17 0.52 0.23 0.52 0.23 1.12 1.125 1.12 1.125 1.25 2.5 1.25 2.5 1.255 2.595 1.255 ;
      POLYGON 2.105 1.15 1.45 1.15 1.45 0.795 1.015 0.795 1.015 0.735 1.45 0.735 1.45 0.36 1.87 0.36 1.87 0.52 1.81 0.52 1.81 0.42 1.51 0.42 1.51 1.09 2.105 1.09 ;
  END
END TLATNCAX4

MACRO TLATNCAX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX6 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.4411 LAYER Metal1 ;
    ANTENNADIFFAREA 2.8394 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.380475 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.4159275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 50.975754 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.14 1.38 4.08 1.38 4.08 0.81 3.73 0.81 3.73 1.38 3.67 1.38 3.67 0.81 3.32 0.81 3.32 1.38 3.26 1.38 3.26 0.35 3.32 0.35 3.32 0.6 3.34 0.6 3.34 0.75 3.67 0.75 3.67 0.35 3.73 0.35 3.73 0.75 4.08 0.75 4.08 0.35 4.14 0.35 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.765 1.335 0.685 1.335 0.685 1.085 0.6 1.085 0.6 0.92 0.68 0.92 0.68 1.005 0.765 1.005 ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.5 1.04 0.42 1.04 0.42 0.895 0.235 0.895 0.235 0.775 0.42 0.775 0.42 0.725 0.5 0.725 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.525 1.65 0.525 1.185 0.585 1.185 0.585 1.65 1.345 1.65 1.345 1.54 1.465 1.54 1.465 1.65 2.195 1.65 2.195 1.51 2.255 1.51 2.255 1.65 2.645 1.65 2.645 1.26 2.705 1.26 2.705 1.65 3.055 1.65 3.055 1.26 3.115 1.26 3.115 1.65 3.465 1.65 3.465 0.91 3.525 0.91 3.525 1.65 3.875 1.65 3.875 0.91 3.935 0.91 3.935 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 3.935 0.06 3.935 0.65 3.875 0.65 3.875 0.06 3.525 0.06 3.525 0.65 3.465 0.65 3.465 0.06 3.065 0.06 3.065 0.47 3.005 0.47 3.005 0.06 2.475 0.06 2.475 0.44 2.355 0.44 2.355 0.38 2.415 0.38 2.415 0.06 1.41 0.06 1.41 0.2 1.35 0.2 1.35 0.06 0.56 0.06 0.56 0.2 0.5 0.2 0.5 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.16 1.1 2.91 1.1 2.91 1.38 2.85 1.38 2.85 1.1 2.5 1.1 2.5 1.38 2.44 1.38 2.44 1.04 3.1 1.04 3.1 0.72 2.845 0.72 2.845 0.56 2.695 0.56 2.695 0.44 2.755 0.44 2.755 0.5 2.905 0.5 2.905 0.66 3.16 0.66 ;
      POLYGON 2.99 0.94 2.355 0.94 2.355 0.76 2.035 0.76 2.035 1.11 1.975 1.11 1.975 0.92 1.345 0.92 1.345 0.86 1.975 0.86 1.975 0.52 2.095 0.52 2.095 0.58 2.035 0.58 2.035 0.7 2.415 0.7 2.415 0.88 2.93 0.88 2.93 0.82 2.99 0.82 ;
      POLYGON 2.68 0.78 2.62 0.78 2.62 0.72 2.535 0.72 2.535 0.6 2.195 0.6 2.195 0.42 1.79 0.42 1.79 0.585 1.73 0.585 1.73 0.76 1.245 0.76 1.245 1.12 1.7 1.12 1.7 1.18 1.185 1.18 1.185 0.7 1.67 0.7 1.67 0.525 1.73 0.525 1.73 0.36 2.255 0.36 2.255 0.54 2.595 0.54 2.595 0.66 2.68 0.66 ;
      POLYGON 2.255 0.92 2.195 0.92 2.195 1.34 0.95 1.34 0.95 1.16 0.865 1.16 0.865 0.53 0.925 0.53 0.925 1.1 1.01 1.1 1.01 1.28 2.135 1.28 2.135 0.86 2.255 0.86 ;
      POLYGON 1.63 0.425 1.57 0.425 1.57 0.43 1.085 0.43 1.085 1 1.025 1 1.025 0.43 0.765 0.43 0.765 0.82 0.705 0.82 0.705 0.625 0.135 0.625 0.135 1.14 0.38 1.14 0.38 1.26 0.32 1.26 0.32 1.2 0.075 1.2 0.075 0.565 0.265 0.565 0.265 0.505 0.325 0.505 0.325 0.565 0.705 0.565 0.705 0.37 1.51 0.37 1.51 0.365 1.63 0.365 ;
  END
END TLATNCAX6

MACRO TLATNCAX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNCAX8 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.618675 LAYER Metal1 ;
    ANTENNADIFFAREA 3.067575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.438075 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.9776865 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 47.498716 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.53 1.395 4.47 1.395 4.47 1.01 4.12 1.01 4.12 1.395 4.06 1.395 4.06 1.01 3.71 1.01 3.71 1.395 3.65 1.395 3.65 1.01 3.3 1.01 3.3 1.395 3.24 1.395 3.24 0.54 3.3 0.54 3.3 0.6 3.34 0.6 3.34 0.95 4.47 0.95 4.47 0.645 3.695 0.645 3.695 0.63 3.62 0.63 3.62 0.57 3.74 0.57 3.74 0.585 4.03 0.585 4.03 0.57 4.15 0.57 4.15 0.585 4.47 0.585 4.47 0.525 4.53 0.525 ;
    END
  END ECK
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.775 1.15 0.535 1.15 0.535 1.07 0.58 1.07 0.58 0.81 0.66 0.81 0.66 1.005 0.775 1.005 ;
    END
  END E
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.435 1.085 0.19 1.085 0.19 1.005 0.355 1.005 0.355 0.75 0.435 0.75 ;
    END
  END CK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.77 0 1.77 0 1.65 0.505 1.65 0.505 1.25 0.565 1.25 0.565 1.65 1.415 1.65 1.415 1.54 1.535 1.54 1.535 1.65 2.185 1.65 2.185 1.51 2.245 1.51 2.245 1.65 2.625 1.65 2.625 1.275 2.685 1.275 2.685 1.65 3.035 1.65 3.035 1.275 3.095 1.275 3.095 1.65 3.445 1.65 3.445 1.11 3.505 1.11 3.505 1.65 3.855 1.65 3.855 1.11 3.915 1.11 3.915 1.65 4.265 1.65 4.265 1.11 4.325 1.11 4.325 1.65 4.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 0.06 4.325 0.06 4.325 0.485 4.265 0.485 4.265 0.06 3.915 0.06 3.915 0.485 3.855 0.485 3.855 0.06 3.505 0.06 3.505 0.485 3.445 0.485 3.445 0.06 3.045 0.06 3.045 0.485 2.985 0.485 2.985 0.06 2.455 0.06 2.455 0.455 2.335 0.455 2.335 0.395 2.395 0.395 2.395 0.06 1.475 0.06 1.475 0.2 1.415 0.2 1.415 0.06 0.51 0.06 0.51 0.49 0.45 0.49 0.45 0.06 0 0.06 0 -0.06 4.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.14 1.115 2.89 1.115 2.89 1.395 2.83 1.395 2.83 1.115 2.48 1.115 2.48 1.395 2.42 1.395 2.42 1.055 3.08 1.055 3.08 0.735 2.825 0.735 2.825 0.575 2.675 0.575 2.675 0.455 2.735 0.455 2.735 0.515 2.885 0.515 2.885 0.675 3.14 0.675 ;
      POLYGON 2.97 0.955 2.355 0.955 2.355 0.775 2.03 0.775 2.03 1.125 1.97 1.125 1.97 0.815 1.415 0.815 1.415 0.755 1.955 0.755 1.955 0.535 2.075 0.535 2.075 0.595 2.015 0.595 2.015 0.715 2.415 0.715 2.415 0.895 2.91 0.895 2.91 0.835 2.97 0.835 ;
      POLYGON 2.66 0.795 2.6 0.795 2.6 0.735 2.515 0.735 2.515 0.615 2.175 0.615 2.175 0.435 1.855 0.435 1.855 0.45 1.795 0.45 1.795 0.655 1.315 0.655 1.315 1.185 1.77 1.185 1.77 1.245 1.255 1.245 1.255 0.655 1.195 0.655 1.195 0.595 1.735 0.595 1.735 0.39 1.795 0.39 1.795 0.375 2.235 0.375 2.235 0.555 2.575 0.555 2.575 0.675 2.66 0.675 ;
      POLYGON 2.25 0.935 2.19 0.935 2.19 1.285 2.085 1.285 2.085 1.405 0.96 1.405 0.96 1.215 0.875 1.215 0.875 0.395 0.935 0.395 0.935 1.155 1.02 1.155 1.02 1.345 2.025 1.345 2.025 1.225 2.13 1.225 2.13 0.875 2.25 0.875 ;
      POLYGON 1.695 0.29 1.635 0.29 1.635 0.36 1.255 0.36 1.255 0.295 1.095 0.295 1.095 0.995 1.035 0.995 1.035 0.295 0.745 0.295 0.745 0.71 0.685 0.71 0.685 0.65 0.09 0.65 0.09 1.185 0.36 1.185 0.36 1.305 0.3 1.305 0.3 1.245 0.03 1.245 0.03 0.59 0.245 0.59 0.245 0.395 0.305 0.395 0.305 0.59 0.685 0.59 0.685 0.235 1.315 0.235 1.315 0.3 1.575 0.3 1.575 0.23 1.695 0.23 ;
  END
END TLATNCAX8

MACRO TLATNSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNSRX1 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.155 LAYER Metal1 ;
    ANTENNADIFFAREA 2.480125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.18495 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.65179775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 87.16950525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 1.33 0.88 1.33 0.88 0.54 0.86 0.54 0.86 0.41 0.94 0.41 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.155 LAYER Metal1 ;
    ANTENNADIFFAREA 2.480125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.18495 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.65179775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 87.16950525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.305 1.29 0.225 1.29 0.225 0.73 0.06 0.73 0.06 0.6 0.225 0.6 0.225 0.54 0.305 0.54 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.245 1.06 4.14 1.06 4.14 1.18 4.06 1.18 4.06 0.98 4.165 0.98 4.165 0.785 4.245 0.785 ;
    END
  END GN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 26.29629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.96 0.905 3.705 0.905 3.705 0.895 3.635 0.895 3.635 0.815 3.705 0.815 3.705 0.36 1.795 0.36 1.795 0.3 3.765 0.3 3.765 0.845 3.96 0.845 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.94 0.92 2.9 0.92 2.9 1.08 2.82 1.08 2.82 0.8 2.86 0.8 2.86 0.62 2.94 0.62 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 0.89 1.28 0.89 1.28 1.11 1.06 1.11 1.06 0.98 1.2 0.98 1.2 0.81 1.34 0.81 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.77 0 1.77 0 1.65 0.475 1.65 0.475 0.9 0.535 0.9 0.535 1.65 1.085 1.65 1.085 1.21 1.145 1.21 1.145 1.65 1.695 1.65 1.695 1.51 1.755 1.51 1.755 1.65 2.1 1.65 2.1 1.51 2.16 1.51 2.16 1.65 2.895 1.65 2.895 1.18 2.955 1.18 2.955 1.65 3.635 1.65 3.635 1.28 3.695 1.28 3.695 1.65 4.11 1.65 4.11 1.28 4.17 1.28 4.17 1.65 4.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 0.06 4.17 0.06 4.17 0.525 4.11 0.525 4.11 0.06 2.915 0.06 2.915 0.2 2.855 0.2 2.855 0.06 1.695 0.06 1.695 0.465 1.85 0.465 1.85 0.525 1.635 0.525 1.635 0.06 1.145 0.06 1.145 0.52 1.085 0.52 1.085 0.06 0.535 0.06 0.535 0.52 0.475 0.52 0.475 0.06 0 0.06 0 -0.06 4.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.405 1.305 4.345 1.305 4.345 0.685 3.925 0.685 3.925 0.745 3.865 0.745 3.865 0.625 4.345 0.625 4.345 0.43 4.405 0.43 ;
      POLYGON 3.9 1.305 3.84 1.305 3.84 1.065 3.475 1.065 3.475 0.71 3.2 0.71 3.2 0.65 3.475 0.65 3.475 0.46 3.605 0.46 3.605 0.52 3.535 0.52 3.535 1.005 3.9 1.005 ;
      POLYGON 3.19 0.525 3.1 0.525 3.1 0.81 3.16 0.81 3.16 1.205 3.1 1.205 3.1 0.87 3.04 0.87 3.04 0.52 2.72 0.52 2.72 0.84 2.355 0.84 2.355 0.78 2.66 0.78 2.66 0.46 3.19 0.46 ;
      POLYGON 2.585 1.205 2.525 1.205 2.525 1 2.195 1 2.195 0.93 1.6 0.93 1.6 0.81 1.66 0.81 1.66 0.87 2.195 0.87 2.195 0.62 2.5 0.62 2.5 0.46 2.56 0.46 2.56 0.68 2.255 0.68 2.255 0.94 2.585 0.94 ;
      RECT 1.835 1.1 2.415 1.18 ;
      POLYGON 2.095 0.71 1.5 0.71 1.5 1.095 1.44 1.095 1.44 0.71 1.1 0.71 1.1 0.82 1.04 0.82 1.04 0.65 1.475 0.65 1.475 0.54 1.535 0.54 1.535 0.65 2.095 0.65 ;
      POLYGON 0.74 1.29 0.68 1.29 0.68 0.79 0.405 0.79 0.405 0.73 0.68 0.73 0.68 0.54 0.74 0.54 ;
  END
END TLATNSRX1

MACRO TLATNSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNSRX2 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.515375 LAYER Metal1 ;
    ANTENNADIFFAREA 3.057325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.279675 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.9939215 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 68.96218825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.14 1.04 4.06 1.04 4.06 0.67 3.985 0.67 3.985 0.51 4.065 0.51 4.065 0.59 4.14 0.59 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.470975 LAYER Metal1 ;
    ANTENNADIFFAREA 3.057325 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.279675 LAYER Metal1 ;
      ANTENNAMAXAREACAR 8.83516575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 68.2810405 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.14 0.98 3.115 0.98 3.115 1.04 3.035 1.04 3.035 0.9 3.06 0.9 3.06 0.51 3.14 0.51 ;
    END
  END QN
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.43 1.04 4.26 1.04 4.26 0.63 4.34 0.63 4.34 0.735 4.43 0.735 ;
    END
  END GN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.66 0.75 2.74 1.25 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 0.92 1.86 0.92 1.86 0.87 1.49 0.87 1.49 0.79 1.94 0.79 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.77777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.755 0.61 1.025 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.43 1.65 0.43 1.285 0.49 1.285 0.49 1.65 1.475 1.65 1.475 1.54 1.595 1.54 1.595 1.65 1.905 1.65 1.905 1.51 1.965 1.51 1.965 1.65 2.58 1.65 2.58 1.51 2.64 1.51 2.64 1.65 2.8 1.65 2.8 1.51 2.86 1.51 2.86 1.65 3.24 1.65 3.24 1.3 3.36 1.3 3.36 1.36 3.3 1.36 3.3 1.65 3.71 1.65 3.71 1.3 3.83 1.3 3.83 1.36 3.77 1.36 3.77 1.65 4.295 1.65 4.295 1.3 4.355 1.3 4.355 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 4.25 0.06 4.25 0.49 4.19 0.49 4.19 0.06 3.77 0.06 3.77 0.49 3.71 0.49 3.71 0.06 3.325 0.06 3.325 0.49 3.265 0.49 3.265 0.06 2.89 0.06 2.89 0.49 2.83 0.49 2.83 0.06 1.835 0.06 1.835 0.19 1.895 0.19 1.895 0.25 1.775 0.25 1.775 0.06 0.41 0.06 0.41 0.435 0.47 0.435 0.47 0.495 0.35 0.495 0.35 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.59 1.2 2.9 1.2 2.9 1.41 2.115 1.41 2.115 1.35 2.84 1.35 2.84 1.14 4.53 1.14 4.53 0.51 4.59 0.51 ;
      POLYGON 3.935 0.85 3.585 0.85 3.585 1.04 3.505 1.04 3.505 0.51 3.585 0.51 3.585 0.77 3.935 0.77 ;
      POLYGON 2.96 0.8 2.9 0.8 2.9 0.65 2.56 0.65 2.56 1.04 2.5 1.04 2.5 0.65 2.445 0.65 2.445 0.33 2.055 0.33 2.055 0.41 1.615 0.41 1.615 0.335 1.5 0.335 1.5 0.275 1.675 0.275 1.675 0.35 1.995 0.35 1.995 0.27 2.505 0.27 2.505 0.59 2.96 0.59 ;
      POLYGON 2.4 0.88 2.32 0.88 2.32 1.25 1.92 1.25 1.92 1.41 1.805 1.41 1.805 1.44 0.985 1.44 0.985 1.04 1.09 1.04 1.09 0.43 1.15 0.43 1.15 1.1 1.045 1.1 1.045 1.38 1.745 1.38 1.745 1.35 1.86 1.35 1.86 1.19 2.26 1.19 2.26 0.82 2.34 0.82 2.34 0.76 2.4 0.76 ;
      POLYGON 2.215 0.69 2.1 0.69 2.1 0.95 2.16 0.95 2.16 1.01 2.04 1.01 2.04 0.69 1.25 0.69 1.25 0.33 0.99 0.33 0.99 0.94 0.93 0.94 0.93 0.655 0.36 0.655 0.36 0.73 0.3 0.73 0.3 0.61 0.315 0.61 0.315 0.595 0.93 0.595 0.93 0.27 1.31 0.27 1.31 0.63 2.155 0.63 2.155 0.43 2.215 0.43 ;
      POLYGON 1.76 1.125 1.33 1.125 1.33 1.28 1.16 1.28 1.16 1.2 1.25 1.2 1.25 1.045 1.76 1.045 ;
      POLYGON 0.83 0.815 0.77 0.815 0.77 1.185 0.285 1.185 0.285 1.31 0.225 1.31 0.225 1.185 0.14 1.185 0.14 0.465 0.175 0.465 0.175 0.405 0.235 0.405 0.235 0.525 0.2 0.525 0.2 1.125 0.71 1.125 0.71 0.755 0.83 0.755 ;
  END
END TLATNSRX2

MACRO TLATNSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNSRX4 0 0 ;
  SIZE 6.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.375475 LAYER Metal1 ;
    ANTENNADIFFAREA 4.29955 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.47835 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.05649625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 54.02947625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.24 1.315 6.18 1.315 6.18 0.92 5.875 0.92 5.875 0.995 5.83 0.995 5.83 1.315 5.77 1.315 5.77 0.935 5.815 0.935 5.815 0.68 5.69 0.68 5.69 0.54 5.75 0.54 5.75 0.62 6.1 0.62 6.1 0.54 6.16 0.54 6.16 0.68 5.94 0.68 5.94 0.86 6.24 0.86 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.375475 LAYER Metal1 ;
    ANTENNADIFFAREA 4.29955 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.47835 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.05649625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 54.02947625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.535 1.315 4.475 1.315 4.475 0.985 4.14 0.985 4.14 1.11 4.125 1.11 4.125 1.315 4.06 1.315 4.06 0.925 4.08 0.925 4.08 0.68 4.05 0.68 4.05 0.54 4.11 0.54 4.11 0.62 4.46 0.62 4.46 0.54 4.52 0.54 4.52 0.68 4.14 0.68 4.14 0.925 4.535 0.925 ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.05178 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.79 0.845 3.765 0.845 3.765 0.895 3.695 0.895 3.695 0.935 3.145 0.935 3.145 0.855 3.085 0.855 3.085 0.795 3.205 0.795 3.205 0.875 3.635 0.875 3.635 0.785 3.79 0.785 ;
    END
  END SN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.66 0.695 1.74 1.195 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 30.18518525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.935 0.36 1.465 0.36 1.465 0.275 0.89 0.275 0.89 0.895 0.635 0.895 0.635 0.875 0.44 0.875 0.44 0.815 0.83 0.815 0.83 0.215 1.525 0.215 1.525 0.3 2.935 0.3 ;
    END
  END RN
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.7 0.34 1.2 ;
    END
  END GN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 1.77 0 1.77 0 1.65 0.3 1.65 0.3 1.51 0.36 1.51 0.36 1.65 0.805 1.65 0.805 1.54 0.925 1.54 0.925 1.65 1.535 1.65 1.535 1.54 1.655 1.54 1.655 1.65 2.5 1.65 2.5 1.34 2.56 1.34 2.56 1.65 3.015 1.65 3.015 1.51 3.075 1.51 3.075 1.65 3.415 1.65 3.415 1.51 3.475 1.51 3.475 1.65 3.86 1.65 3.86 1.195 3.92 1.195 3.92 1.65 4.27 1.65 4.27 1.085 4.33 1.085 4.33 1.65 4.68 1.65 4.68 0.925 4.74 0.925 4.74 1.65 5.09 1.65 5.09 0.925 5.15 0.925 5.15 1.65 5.5 1.65 5.5 0.94 5.56 0.94 5.56 1.65 5.975 1.65 5.975 1.02 6.035 1.02 6.035 1.65 6.385 1.65 6.385 0.925 6.445 0.925 6.445 1.65 6.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.6 0.06 6.365 0.06 6.365 0.52 6.305 0.52 6.305 0.06 5.955 0.06 5.955 0.52 5.895 0.52 5.895 0.06 5.545 0.06 5.545 0.52 5.485 0.52 5.485 0.06 5.135 0.06 5.135 0.52 5.075 0.52 5.075 0.06 4.725 0.06 4.725 0.52 4.665 0.52 4.665 0.06 4.315 0.06 4.315 0.52 4.255 0.52 4.255 0.06 3.885 0.06 3.885 0.52 3.825 0.52 3.825 0.06 3.11 0.06 3.11 0.52 3.05 0.52 3.05 0.06 1.845 0.06 1.845 0.2 1.785 0.2 1.785 0.06 1.685 0.06 1.685 0.2 1.625 0.2 1.625 0.06 0.455 0.06 0.455 0.44 0.395 0.44 0.395 0.06 0 0.06 0 -0.06 6.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.715 0.84 5.31 0.84 5.31 0.94 5.355 0.94 5.355 1.315 5.295 1.315 5.295 1 5.25 1 5.25 0.825 4.945 0.825 4.945 1.315 4.885 1.315 4.885 0.66 4.87 0.66 4.87 0.54 4.93 0.54 4.93 0.6 4.945 0.6 4.945 0.765 5.28 0.765 5.28 0.54 5.34 0.54 5.34 0.78 5.715 0.78 ;
      POLYGON 3.95 1.095 3.64 1.095 3.64 1.155 3.58 1.155 3.58 1.095 3.24 1.095 3.24 1.155 3.18 1.155 3.18 1.095 2.925 1.095 2.925 0.965 2.71 0.965 2.71 0.905 2.985 0.905 2.985 1.035 3.89 1.035 3.89 0.685 3.465 0.685 3.465 0.485 3.525 0.485 3.525 0.625 3.95 0.625 ;
      POLYGON 3.365 0.775 3.305 0.775 3.305 0.695 2.61 0.695 2.61 1.06 2.075 1.06 2.075 1.12 2.06 1.12 2.06 1.18 2 1.18 2 1.06 2.015 1.06 2.015 1 2.55 1 2.55 0.695 2.33 0.695 2.33 0.58 2.295 0.58 2.295 0.46 2.355 0.46 2.355 0.52 2.39 0.52 2.39 0.635 3.365 0.635 ;
      RECT 2.175 1.16 2.825 1.24 ;
      POLYGON 2.45 0.9 1.9 0.9 1.9 1.355 1.5 1.355 1.5 1.375 0.99 1.375 0.99 1.055 0.66 1.055 0.66 1.245 0.6 1.245 0.6 0.995 0.99 0.995 0.99 0.375 1.11 0.375 1.11 0.435 1.05 0.435 1.05 1.315 1.44 1.315 1.44 0.82 1.56 0.82 1.56 0.88 1.5 0.88 1.5 1.295 1.84 1.295 1.84 0.84 2.45 0.84 ;
      POLYGON 2.23 0.74 2.11 0.74 2.11 0.595 1.34 0.595 1.34 1.215 1.22 1.215 1.22 1.155 1.28 1.155 1.28 0.535 1.3 0.535 1.3 0.515 1.42 0.515 1.42 0.535 2.17 0.535 2.17 0.68 2.23 0.68 ;
      POLYGON 0.73 0.6 0.13 0.6 0.13 1.34 0.07 1.34 0.07 0.54 0.19 0.54 0.19 0.345 0.25 0.345 0.25 0.54 0.73 0.54 ;
  END
END TLATNSRX4

MACRO TLATNSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNSRXL 0 0 ;
  SIZE 4.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.14115 LAYER Metal1 ;
    ANTENNADIFFAREA 2.381075 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1458 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.685528 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 107.22222225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.055 0.625 0.94 0.625 0.94 1.03 1.055 1.03 1.055 1.175 0.975 1.175 0.975 1.11 0.86 1.11 0.86 0.545 0.975 0.545 0.975 0.505 1.055 0.505 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.14115 LAYER Metal1 ;
    ANTENNADIFFAREA 2.381075 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1458 LAYER Metal1 ;
      ANTENNAMAXAREACAR 14.685528 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 107.22222225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.325 1.02 0.245 1.02 0.245 0.73 0.06 0.73 0.06 0.6 0.245 0.6 0.245 0.54 0.325 0.54 ;
    END
  END Q
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.41 1.11 4.34 1.11 4.34 1.26 4.26 1.26 4.26 0.83 4.41 0.83 ;
    END
  END GN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 27.45370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.16 0.92 3.66 0.92 3.66 0.79 3.73 0.79 3.73 0.405 1.84 0.405 1.84 0.345 3.79 0.345 3.79 0.86 4.16 0.86 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.18 0.92 3.025 0.92 3.025 1.01 2.945 1.01 2.945 0.665 3.18 0.665 ;
    END
  END D
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.365 1.275 1.175 1.275 1.175 1.195 1.285 1.195 1.285 0.885 1.365 0.885 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 1.77 0 1.77 0 1.65 0.525 1.65 0.525 1.285 0.585 1.285 0.585 1.65 1.23 1.65 1.23 1.51 1.29 1.51 1.29 1.65 1.745 1.65 1.745 1.51 1.805 1.51 1.805 1.65 2.145 1.65 2.145 1.265 2.205 1.265 2.205 1.65 2.99 1.65 2.99 1.11 3.05 1.11 3.05 1.65 3.72 1.65 3.72 1.36 3.78 1.36 3.78 1.65 4.21 1.65 4.21 1.36 4.27 1.36 4.27 1.65 4.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.6 0.06 4.27 0.06 4.27 0.57 4.21 0.57 4.21 0.06 3.08 0.06 3.08 0.2 3.02 0.2 3.02 0.06 1.74 0.06 1.74 0.54 1.895 0.54 1.895 0.6 1.68 0.6 1.68 0.06 1.26 0.06 1.26 0.62 1.2 0.62 1.2 0.06 0.555 0.06 0.555 0.635 0.495 0.635 0.495 0.06 0 0.06 0 -0.06 4.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.57 1.325 4.5 1.325 4.5 1.385 4.44 1.385 4.44 1.265 4.51 1.265 4.51 0.73 3.89 0.73 3.89 0.67 4.47 0.67 4.47 0.475 4.57 0.475 ;
      POLYGON 4.045 1.385 3.985 1.385 3.985 1.26 3.5 1.26 3.5 0.79 3.44 0.79 3.44 0.73 3.5 0.73 3.5 0.505 3.63 0.505 3.63 0.565 3.56 0.565 3.56 1.2 4.045 1.2 ;
      POLYGON 3.4 0.63 3.34 0.63 3.34 1.135 3.28 1.135 3.28 0.565 2.845 0.565 2.845 0.815 2.48 0.815 2.48 0.825 2.36 0.825 2.36 0.765 2.42 0.765 2.42 0.755 2.785 0.755 2.785 0.505 3.4 0.505 ;
      POLYGON 2.685 0.655 2.26 0.655 2.26 0.925 2.58 0.925 2.58 1.135 2.52 1.135 2.52 0.985 1.625 0.985 1.625 0.925 2.2 0.925 2.2 0.595 2.625 0.595 2.625 0.535 2.685 0.535 ;
      RECT 1.88 1.085 2.405 1.165 ;
      POLYGON 2.1 0.825 2.04 0.825 2.04 0.785 1.525 0.785 1.525 1.175 1.465 1.175 1.465 0.785 1.095 0.785 1.095 0.725 1.52 0.725 1.52 0.525 1.58 0.525 1.58 0.725 2.04 0.725 2.04 0.705 2.1 0.705 ;
      POLYGON 0.76 1.02 0.68 1.02 0.68 0.815 0.425 0.815 0.425 0.735 0.68 0.735 0.68 0.54 0.76 0.54 ;
  END
END TLATNSRXL

MACRO TLATNTSCAX12
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX12 0 0 ;
  SIZE 6.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.72865 LAYER Metal1 ;
    ANTENNADIFFAREA 4.377425 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.62055 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.0086215 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 48.18950925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.935 0.85 5.89 0.85 5.89 0.95 5.935 0.95 5.935 1.42 5.875 1.42 5.875 1.01 5.83 1.01 5.83 0.85 5.525 0.85 5.525 1.42 5.465 1.42 5.465 0.85 5.115 0.85 5.115 1.42 5.055 1.42 5.055 0.85 4.705 0.85 4.705 1.42 4.645 1.42 4.645 0.85 4.34 0.85 4.34 0.92 4.3 0.92 4.3 0.925 4.295 0.925 4.295 1.42 4.235 1.42 4.235 0.87 4.26 0.87 4.26 0.66 4.235 0.66 4.235 0.35 4.295 0.35 4.295 0.605 4.32 0.605 4.32 0.79 4.645 0.79 4.645 0.35 4.705 0.35 4.705 0.79 5.055 0.79 5.055 0.35 5.115 0.35 5.115 0.79 5.465 0.79 5.465 0.35 5.525 0.35 5.525 0.79 5.875 0.79 5.875 0.35 5.935 0.35 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.745 0.945 0.665 0.945 0.665 0.73 0.66 0.73 0.66 0.45 0.745 0.45 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.64814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.45 0.54 0.945 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 12.037037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.205 0.56 0.14 0.56 0.14 0.945 0.06 0.945 0.06 0.44 0.205 0.44 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 1.77 0 1.77 0 1.65 0.525 1.65 0.525 1.21 0.585 1.21 0.585 1.65 1.765 1.65 1.765 1.55 1.705 1.55 1.705 1.49 1.825 1.49 1.825 1.65 2.565 1.65 2.565 1.03 2.625 1.03 2.625 1.65 3.045 1.65 3.045 1.3 3.105 1.3 3.105 1.65 3.455 1.65 3.455 1.3 3.515 1.3 3.515 1.65 3.9 1.65 3.9 1.33 4.02 1.33 4.02 1.39 3.96 1.39 3.96 1.65 4.44 1.65 4.44 0.95 4.5 0.95 4.5 1.65 4.85 1.65 4.85 0.95 4.91 0.95 4.91 1.65 5.26 1.65 5.26 0.95 5.32 0.95 5.32 1.65 5.67 1.65 5.67 0.95 5.73 0.95 5.73 1.65 6.08 1.65 6.08 0.95 6.14 0.95 6.14 1.65 6.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 6.4 0.06 6.14 0.06 6.14 0.66 6.08 0.66 6.08 0.06 5.73 0.06 5.73 0.66 5.67 0.66 5.67 0.06 5.32 0.06 5.32 0.66 5.26 0.66 5.26 0.06 4.91 0.06 4.91 0.66 4.85 0.66 4.85 0.06 4.5 0.06 4.5 0.66 4.44 0.66 4.44 0.06 4.09 0.06 4.09 0.47 4.03 0.47 4.03 0.06 3.385 0.06 3.385 0.41 3.445 0.41 3.445 0.47 3.325 0.47 3.325 0.06 2.73 0.06 2.73 0.43 2.67 0.43 2.67 0.06 1.705 0.06 1.705 0.25 1.765 0.25 1.765 0.31 1.645 0.31 1.645 0.06 0.585 0.06 0.585 0.35 0.525 0.35 0.525 0.06 0.155 0.06 0.155 0.35 0.095 0.35 0.095 0.06 0 0.06 0 -0.06 6.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.16 0.795 4.015 0.795 4.015 1.11 3.785 1.11 3.785 1.42 3.725 1.42 3.725 1.11 3.31 1.11 3.31 1.42 3.25 1.42 3.25 1.11 2.9 1.11 2.9 1.37 2.84 1.37 2.84 1.05 3.955 1.05 3.955 0.63 3.085 0.63 3.085 0.61 3.015 0.61 3.015 0.55 3.135 0.55 3.135 0.57 3.83 0.57 3.83 0.51 3.89 0.51 3.89 0.57 4.015 0.57 4.015 0.735 4.16 0.735 ;
      POLYGON 3.855 0.79 2.855 0.79 2.855 0.59 2.51 0.59 2.51 0.42 2.145 0.42 2.145 0.595 2.085 0.595 2.085 0.855 1.74 0.855 1.74 1.115 2.145 1.115 2.145 1.21 2.205 1.21 2.205 1.27 2.085 1.27 2.085 1.175 1.68 1.175 1.68 0.92 1.62 0.92 1.62 0.795 2.025 0.795 2.025 0.535 2.085 0.535 2.085 0.36 2.57 0.36 2.57 0.53 2.915 0.53 2.915 0.73 3.855 0.73 ;
      POLYGON 3.37 0.95 2.695 0.95 2.695 0.75 2.305 0.75 2.305 1.1 2.245 1.1 2.245 1.015 1.84 1.015 1.84 0.955 2.245 0.955 2.245 0.69 2.35 0.69 2.35 0.52 2.41 0.52 2.41 0.69 2.755 0.69 2.755 0.89 3.37 0.89 ;
      POLYGON 2.59 0.91 2.465 0.91 2.465 1.43 1.925 1.43 1.925 1.335 1.455 1.335 1.455 1.395 1.395 1.395 1.395 1.335 1.3 1.335 1.3 0.63 1.24 0.63 1.24 0.57 1.36 0.57 1.36 1.275 1.985 1.275 1.985 1.37 2.405 1.37 2.405 0.85 2.59 0.85 ;
      POLYGON 1.985 0.435 1.925 0.435 1.925 0.47 1.52 0.47 1.52 1.14 1.46 1.14 1.46 0.47 1.22 0.47 1.22 0.315 0.905 0.315 0.905 1.235 0.845 1.235 0.845 0.375 0.82 0.375 0.82 0.255 1.28 0.255 1.28 0.41 1.865 0.41 1.865 0.375 1.985 0.375 ;
      POLYGON 1.2 1.395 0.685 1.395 0.685 1.11 0.275 1.11 0.275 1.235 0.215 1.235 0.215 1.05 0.3 1.05 0.3 0.255 0.36 0.255 0.36 1.05 0.745 1.05 0.745 1.335 1.08 1.335 1.08 0.63 1.02 0.63 1.02 0.57 1.14 0.57 1.14 1.275 1.2 1.275 ;
  END
END TLATNTSCAX12

MACRO TLATNTSCAX16
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX16 0 0 ;
  SIZE 7.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.395 LAYER Metal1 ;
    ANTENNADIFFAREA 5.224225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.81135 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.41689775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 43.1798855 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.18 1.405 7.12 1.405 7.12 0.875 6.77 0.875 6.77 1.405 6.71 1.405 6.71 0.875 6.36 0.875 6.36 1.405 6.3 1.405 6.3 0.875 5.95 0.875 5.95 1.405 5.89 1.405 5.89 0.875 5.54 0.875 5.54 1.405 5.48 1.405 5.48 0.875 5.13 0.875 5.13 1.405 5.07 1.405 5.07 0.875 4.74 0.875 4.74 0.92 4.72 0.92 4.72 1.405 4.66 1.405 4.66 0.62 4.615 0.62 4.615 0.5 4.675 0.5 4.675 0.56 4.72 0.56 4.72 0.79 4.74 0.79 4.74 0.815 5.435 0.815 5.435 0.645 5.07 0.645 5.07 0.63 4.995 0.63 4.995 0.57 5.115 0.57 5.115 0.585 5.435 0.585 5.435 0.525 5.495 0.525 5.495 0.815 6.255 0.815 6.255 0.645 5.89 0.645 5.89 0.63 5.815 0.63 5.815 0.57 5.935 0.57 5.935 0.585 6.255 0.585 6.255 0.525 6.315 0.525 6.315 0.815 7.075 0.815 7.075 0.645 6.71 0.645 6.71 0.63 6.635 0.63 6.635 0.57 6.755 0.57 6.755 0.585 7.075 0.585 7.075 0.525 7.135 0.525 7.135 0.815 7.18 0.815 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.45 0.74 0.95 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.45 0.54 0.95 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.27777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.145 0.95 0.06 0.95 0.06 0.48 0.14 0.48 0.14 0.83 0.145 0.83 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.6 1.77 0 1.77 0 1.65 0.46 1.65 0.46 1.27 0.4 1.27 0.4 1.21 0.52 1.21 0.52 1.65 1.665 1.65 1.665 1.305 1.785 1.305 1.785 1.365 1.725 1.365 1.725 1.65 2.275 1.65 2.275 1.51 2.335 1.51 2.335 1.65 2.795 1.65 2.795 1.095 2.855 1.095 2.855 1.65 3.225 1.65 3.225 1.285 3.285 1.285 3.285 1.65 3.635 1.65 3.635 1.285 3.695 1.285 3.695 1.65 4.045 1.65 4.045 1.285 4.105 1.285 4.105 1.65 4.455 1.65 4.455 1.285 4.515 1.285 4.515 1.65 4.865 1.65 4.865 0.975 4.925 0.975 4.925 1.65 5.275 1.65 5.275 0.975 5.335 0.975 5.335 1.65 5.685 1.65 5.685 0.975 5.745 0.975 5.745 1.65 6.095 1.65 6.095 0.975 6.155 0.975 6.155 1.65 6.505 1.65 6.505 0.975 6.565 0.975 6.565 1.65 6.915 1.65 6.915 0.975 6.975 0.975 6.975 1.65 7.325 1.65 7.325 0.96 7.385 0.96 7.385 1.65 7.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.6 0.06 7.34 0.06 7.34 0.485 7.28 0.485 7.28 0.06 6.93 0.06 6.93 0.485 6.87 0.485 6.87 0.06 6.52 0.06 6.52 0.485 6.46 0.485 6.46 0.06 6.11 0.06 6.11 0.485 6.05 0.485 6.05 0.06 5.7 0.06 5.7 0.485 5.64 0.485 5.64 0.06 5.29 0.06 5.29 0.485 5.23 0.485 5.23 0.06 4.88 0.06 4.88 0.485 4.82 0.485 4.82 0.06 4.47 0.06 4.47 0.485 4.41 0.485 4.41 0.06 3.765 0.06 3.765 0.395 3.825 0.395 3.825 0.455 3.705 0.455 3.705 0.06 3.125 0.06 3.125 0.575 3.065 0.575 3.065 0.06 2.57 0.06 2.57 0.17 2.45 0.17 2.45 0.06 1.975 0.06 1.975 0.25 1.855 0.25 1.855 0.19 1.915 0.19 1.915 0.06 0.585 0.06 0.585 0.35 0.525 0.35 0.525 0.06 0.155 0.06 0.155 0.35 0.095 0.35 0.095 0.06 0 0.06 0 -0.06 7.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.56 1.095 4.31 1.095 4.31 1.405 4.25 1.405 4.25 1.095 3.9 1.095 3.9 1.405 3.84 1.405 3.84 1.095 3.49 1.095 3.49 1.405 3.43 1.405 3.43 1.095 3.08 1.095 3.08 1.405 3.02 1.405 3.02 1.035 4.5 1.035 4.5 0.775 4.25 0.775 4.25 0.615 3.555 0.615 3.555 0.595 3.345 0.595 3.345 0.535 3.605 0.535 3.605 0.555 4.045 0.555 4.045 0.495 4.105 0.495 4.105 0.555 4.31 0.555 4.31 0.715 4.56 0.715 ;
      POLYGON 4.4 0.935 2.695 0.935 2.695 1.185 2.57 1.185 2.57 1.405 2.51 1.405 2.51 1.125 2.635 1.125 2.635 0.865 1.78 0.865 1.78 0.725 1.84 0.725 1.84 0.805 2.685 0.805 2.685 0.57 2.805 0.57 2.805 0.63 2.745 0.63 2.745 0.875 4.4 0.875 ;
      POLYGON 4.06 0.775 2.905 0.775 2.905 0.47 2.355 0.47 2.355 0.565 2.295 0.565 2.295 0.625 1.68 0.625 1.68 0.985 2.105 0.985 2.105 1.055 2.165 1.055 2.165 1.115 2.045 1.115 2.045 1.045 1.62 1.045 1.62 0.565 2.235 0.565 2.235 0.505 2.295 0.505 2.295 0.41 2.965 0.41 2.965 0.715 4.06 0.715 ;
      POLYGON 2.535 1.025 2.325 1.025 2.325 1.275 1.885 1.275 1.885 1.205 1.61 1.205 1.61 1.21 1.445 1.21 1.445 1.3 1.385 1.3 1.385 1.21 1.3 1.21 1.3 0.525 1.36 0.525 1.36 1.15 1.575 1.15 1.575 1.145 1.945 1.145 1.945 1.215 2.265 1.215 2.265 0.965 2.535 0.965 ;
      POLYGON 2.195 0.405 2.135 0.405 2.135 0.41 1.695 0.41 1.695 0.29 1.52 0.29 1.52 1.05 1.46 1.05 1.46 0.29 0.9 0.29 0.9 1.175 0.78 1.175 0.78 1.115 0.84 1.115 0.84 0.35 0.735 0.35 0.735 0.23 1.205 0.23 1.205 0.19 1.325 0.19 1.325 0.23 1.755 0.23 1.755 0.35 2.075 0.35 2.075 0.345 2.195 0.345 ;
      POLYGON 1.155 1.395 1.095 1.395 1.095 1.335 0.62 1.335 0.62 1.11 0.18 1.11 0.18 1.205 0.12 1.205 0.12 1.05 0.3 1.05 0.3 0.255 0.36 0.255 0.36 1.05 0.68 1.05 0.68 1.275 1.095 1.275 1.095 0.525 1.155 0.525 ;
  END
END TLATNTSCAX16

MACRO TLATNTSCAX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX2 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.16 LAYER Metal1 ;
    ANTENNADIFFAREA 2.05005 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1719 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.565445 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 99.21465975 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.36 0.53 3.34 0.53 3.34 1.29 3.26 1.29 3.26 0.41 3.36 0.41 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.45 0.74 0.95 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.45 0.54 0.95 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.79629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.06 0.47 0.14 0.865 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 1.77 0 1.77 0 1.65 0.52 1.65 0.52 1.21 0.58 1.21 0.58 1.65 1.64 1.65 1.64 1.49 1.76 1.49 1.76 1.55 1.7 1.55 1.7 1.65 2.61 1.65 2.61 1.01 2.67 1.01 2.67 1.65 3.055 1.65 3.055 1.01 3.115 1.01 3.115 1.65 3.465 1.65 3.465 0.9 3.525 0.9 3.525 1.65 3.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 0.06 3.565 0.06 3.565 0.52 3.505 0.52 3.505 0.06 3.125 0.06 3.125 0.2 3.065 0.2 3.065 0.06 2.73 0.06 2.73 0.2 2.67 0.2 2.67 0.06 1.79 0.06 1.79 0.53 1.89 0.53 1.89 0.59 1.73 0.59 1.73 0.06 0.58 0.06 0.58 0.35 0.52 0.35 0.52 0.06 0.155 0.06 0.155 0.35 0.095 0.35 0.095 0.06 0 0.06 0 -0.06 3.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.16 0.835 2.955 0.835 2.955 0.995 2.895 0.995 2.895 1.035 2.815 1.035 2.815 0.915 2.875 0.915 2.875 0.755 2.945 0.755 2.945 0.65 2.905 0.65 2.905 0.57 3.025 0.57 3.025 0.755 3.16 0.755 ;
      POLYGON 2.95 0.435 2.21 0.435 2.21 0.91 1.645 0.91 1.645 1.17 2.08 1.17 2.08 1.27 2.14 1.27 2.14 1.33 2.02 1.33 2.02 1.23 1.585 1.23 1.585 0.91 1.525 0.91 1.525 0.85 2.15 0.85 2.15 0.375 2.95 0.375 ;
      POLYGON 2.775 0.8 2.41 0.8 2.41 1.01 2.435 1.01 2.435 1.13 2.375 1.13 2.375 1.07 1.745 1.07 1.745 1.01 2.35 1.01 2.35 0.54 2.41 0.54 2.41 0.74 2.775 0.74 ;
      POLYGON 2.51 1.49 1.86 1.49 1.86 1.39 1.33 1.39 1.33 1.23 1.205 1.23 1.205 0.525 1.265 0.525 1.265 1.17 1.39 1.17 1.39 1.33 1.92 1.33 1.92 1.43 2.45 1.43 2.45 1.23 2.51 1.23 ;
      POLYGON 2.05 0.75 1.57 0.75 1.57 0.29 1.425 0.29 1.425 1.01 1.485 1.01 1.485 1.07 1.365 1.07 1.365 0.29 0.9 0.29 0.9 1.235 0.84 1.235 0.84 0.35 0.735 0.35 0.735 0.23 1.63 0.23 1.63 0.69 1.99 0.69 1.99 0.42 1.89 0.42 1.89 0.36 2.05 0.36 ;
      POLYGON 1.105 1.455 1.045 1.455 1.045 1.395 0.68 1.395 0.68 1.11 0.27 1.11 0.27 1.235 0.21 1.235 0.21 1.05 0.3 1.05 0.3 0.255 0.36 0.255 0.36 1.05 0.74 1.05 0.74 1.335 1.045 1.335 1.045 0.645 1 0.645 1 0.525 1.06 0.525 1.06 0.585 1.105 0.585 ;
  END
END TLATNTSCAX2

MACRO TLATNTSCAX20
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX20 0 0 ;
  SIZE 8.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.281175 LAYER Metal1 ;
    ANTENNADIFFAREA 6.1327 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 1.0008 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.2769535 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 42.26918475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.6 0.66 8.555 0.66 8.555 0.76 8.6 0.76 8.6 1.355 8.54 1.355 8.54 0.82 8.19 0.82 8.19 1.36 8.13 1.36 8.13 0.82 7.78 0.82 7.78 1.36 7.72 1.36 7.72 0.82 7.37 0.82 7.37 1.36 7.31 1.36 7.31 0.82 6.96 0.82 6.96 1.36 6.9 1.36 6.9 0.82 6.55 0.82 6.55 1.36 6.49 1.36 6.49 0.82 6.14 0.82 6.14 1.36 6.08 1.36 6.08 0.82 5.73 0.82 5.73 1.36 5.67 1.36 5.67 0.82 5.34 0.82 5.34 1.36 5.26 1.36 5.26 0.355 5.32 0.355 5.32 0.76 5.67 0.76 5.67 0.355 5.73 0.355 5.73 0.76 6.035 0.76 6.035 0.6 6.08 0.6 6.08 0.355 6.14 0.355 6.14 0.66 6.095 0.66 6.095 0.76 6.49 0.76 6.49 0.355 6.55 0.355 6.55 0.76 6.9 0.76 6.9 0.355 6.96 0.355 6.96 0.76 7.31 0.76 7.31 0.355 7.37 0.355 7.37 0.76 7.72 0.76 7.72 0.355 7.78 0.355 7.78 0.76 8.13 0.76 8.13 0.355 8.19 0.355 8.19 0.76 8.495 0.76 8.495 0.6 8.54 0.6 8.54 0.355 8.6 0.355 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.05 0.895 0.695 0.895 0.695 0.815 0.74 0.815 0.74 0.67 0.965 0.67 0.965 0.815 1.05 0.815 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.595 0.87 0.54 0.87 0.54 0.955 0.46 0.955 0.46 0.79 0.515 0.79 0.515 0.51 0.595 0.51 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.2 1.06 0.14 1.06 0.14 1.14 0.06 1.14 0.06 0.98 0.12 0.98 0.12 0.7 0.2 0.7 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.8 1.77 0 1.77 0 1.65 0.64 1.65 0.64 0.995 0.7 0.995 0.7 1.65 2.01 1.65 2.01 1.345 2.07 1.345 2.07 1.65 2.395 1.65 2.395 1.27 2.515 1.27 2.515 1.33 2.455 1.33 2.455 1.65 2.945 1.65 2.945 1.27 3.065 1.27 3.065 1.33 3.005 1.33 3.005 1.65 3.385 1.65 3.385 1.13 3.445 1.13 3.445 1.65 3.795 1.65 3.795 1.13 3.855 1.13 3.855 1.65 4.205 1.65 4.205 1.13 4.265 1.13 4.265 1.65 4.615 1.65 4.615 1.13 4.675 1.13 4.675 1.65 5.025 1.65 5.025 1.13 5.085 1.13 5.085 1.65 5.465 1.65 5.465 0.92 5.525 0.92 5.525 1.65 5.875 1.65 5.875 0.92 5.935 0.92 5.935 1.65 6.285 1.65 6.285 0.92 6.345 0.92 6.345 1.65 6.695 1.65 6.695 0.92 6.755 0.92 6.755 1.65 7.105 1.65 7.105 0.92 7.165 0.92 7.165 1.65 7.515 1.65 7.515 0.92 7.575 0.92 7.575 1.65 7.925 1.65 7.925 0.92 7.985 0.92 7.985 1.65 8.335 1.65 8.335 0.92 8.395 0.92 8.395 1.65 8.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 8.8 0.06 8.395 0.06 8.395 0.66 8.335 0.66 8.335 0.06 7.985 0.06 7.985 0.66 7.925 0.66 7.925 0.06 7.575 0.06 7.575 0.66 7.515 0.66 7.515 0.06 7.165 0.06 7.165 0.66 7.105 0.66 7.105 0.06 6.755 0.06 6.755 0.66 6.695 0.66 6.695 0.06 6.345 0.06 6.345 0.66 6.285 0.66 6.285 0.06 5.935 0.06 5.935 0.66 5.875 0.66 5.875 0.06 5.525 0.06 5.525 0.66 5.465 0.66 5.465 0.06 5.115 0.06 5.115 0.475 5.055 0.475 5.055 0.06 4.445 0.06 4.445 0.28 4.505 0.28 4.505 0.34 4.385 0.34 4.385 0.06 3.825 0.06 3.825 0.28 3.885 0.28 3.885 0.34 3.765 0.34 3.765 0.06 3.17 0.06 3.17 0.37 3.11 0.37 3.11 0.06 2.76 0.06 2.76 0.37 2.7 0.37 2.7 0.06 2 0.06 2 0.25 2.06 0.25 2.06 0.31 1.94 0.31 1.94 0.06 0.73 0.06 0.73 0.17 0.61 0.17 0.61 0.06 0.2 0.06 0.2 0.6 0.14 0.6 0.14 0.06 0 0.06 0 -0.06 8.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 5.16 0.79 5.1 0.79 5.1 1.03 4.88 1.03 4.88 1.36 4.82 1.36 4.82 1.03 4.47 1.03 4.47 1.36 4.41 1.36 4.41 1.03 4.06 1.03 4.06 1.36 4 1.36 4 1.03 3.65 1.03 3.65 1.36 3.59 1.36 3.59 1.03 3.24 1.03 3.24 1.36 3.18 1.36 3.18 0.97 5.04 0.97 5.04 0.635 4.725 0.635 4.725 0.5 3.525 0.5 3.525 0.48 3.455 0.48 3.455 0.42 3.575 0.42 3.575 0.44 4.075 0.44 4.075 0.42 4.195 0.42 4.195 0.44 4.725 0.44 4.725 0.38 4.785 0.38 4.785 0.575 5.1 0.575 5.1 0.73 5.16 0.73 ;
      POLYGON 4.94 0.865 3.08 0.865 3.08 1.17 2.47 1.17 2.47 1.01 1.79 1.01 1.79 0.57 2.32 0.57 2.32 0.47 2.44 0.47 2.44 0.53 2.38 0.53 2.38 0.63 1.85 0.63 1.85 0.95 2.53 0.95 2.53 1.11 3.02 1.11 3.02 0.805 4.94 0.805 ;
      POLYGON 4.57 0.67 2.92 0.67 2.92 0.85 2.69 0.85 2.69 0.95 2.75 0.95 2.75 1.01 2.63 1.01 2.63 0.85 1.95 0.85 1.95 0.73 2.01 0.73 2.01 0.79 2.86 0.79 2.86 0.45 2.905 0.45 2.905 0.39 2.965 0.39 2.965 0.51 2.92 0.51 2.92 0.61 4.57 0.61 ;
      POLYGON 2.76 0.69 2.49 0.69 2.49 0.63 2.7 0.63 2.7 0.53 2.54 0.53 2.54 0.37 2.22 0.37 2.22 0.47 1.69 0.47 1.69 1.11 1.75 1.11 1.75 1.17 1.63 1.17 1.63 0.35 1.69 0.35 1.69 0.41 2.16 0.41 2.16 0.31 2.6 0.31 2.6 0.47 2.76 0.47 ;
      POLYGON 2.29 1.245 1.91 1.245 1.91 1.33 1.825 1.33 1.825 1.45 1.705 1.45 1.705 1.33 1.435 1.33 1.435 1.265 0.845 1.265 0.845 0.995 1.15 0.995 1.15 0.57 0.87 0.57 0.87 0.51 1.21 0.51 1.21 1.055 0.905 1.055 0.905 1.205 1.47 1.205 1.47 0.58 1.53 0.58 1.53 1.27 1.85 1.27 1.85 1.185 2.29 1.185 ;
      POLYGON 1.48 0.47 1.37 0.47 1.37 1.105 1.31 1.105 1.31 0.41 0.405 0.41 0.405 0.6 0.36 0.6 0.36 1.02 0.3 1.02 0.3 0.54 0.345 0.54 0.345 0.35 1.48 0.35 ;
  END
END TLATNTSCAX20

MACRO TLATNTSCAX3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX3 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.2865 LAYER Metal1 ;
    ANTENNADIFFAREA 2.33575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.22725 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.06160625 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 80.46204625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.93 0.66 3.54 0.66 3.54 0.73 3.52 0.73 3.52 0.9 3.885 0.9 3.885 1.29 3.825 1.29 3.825 0.96 3.475 0.96 3.475 1.29 3.415 1.29 3.415 0.9 3.46 0.9 3.46 0.52 3.52 0.52 3.52 0.6 3.87 0.6 3.87 0.52 3.93 0.52 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.45 0.765 0.925 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 0.73 0.515 0.73 0.515 0.925 0.435 0.925 0.435 0.6 0.46 0.6 0.46 0.45 0.54 0.45 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.64814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.16 0.605 0.14 0.605 0.14 0.95 0.06 0.95 0.06 0.475 0.14 0.475 0.14 0.485 0.16 0.485 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 0 1.77 0 1.65 0.5 1.65 0.5 1.185 0.56 1.185 0.56 1.65 1.755 1.65 1.755 1.49 1.875 1.49 1.875 1.55 1.815 1.55 1.815 1.65 2.73 1.65 2.73 0.995 2.79 0.995 2.79 1.65 3.14 1.65 3.14 1.09 3.2 1.09 3.2 1.65 3.62 1.65 3.62 1.06 3.68 1.06 3.68 1.65 4 1.65 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.725 0.06 3.725 0.5 3.665 0.5 3.665 0.06 3.285 0.06 3.285 0.2 3.225 0.2 3.225 0.06 2.79 0.06 2.79 0.17 2.67 0.17 2.67 0.06 1.905 0.06 1.905 0.53 2.005 0.53 2.005 0.59 1.845 0.59 1.845 0.06 0.56 0.06 0.56 0.35 0.5 0.35 0.5 0.06 0.13 0.06 0.13 0.35 0.07 0.35 0.07 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.36 0.8 3.185 0.8 3.185 0.99 2.995 0.99 2.995 1.29 2.935 1.29 2.935 0.93 3.125 0.93 3.125 0.61 3.095 0.61 3.095 0.49 3.155 0.49 3.155 0.55 3.185 0.55 3.185 0.74 3.36 0.74 ;
      POLYGON 3.025 0.83 2.935 0.83 2.935 0.47 2.325 0.47 2.325 0.91 1.76 0.91 1.76 1.17 2.195 1.17 2.195 1.245 2.255 1.245 2.255 1.305 2.135 1.305 2.135 1.23 1.7 1.23 1.7 0.91 1.64 0.91 1.64 0.85 2.265 0.85 2.265 0.41 2.995 0.41 2.995 0.71 3.025 0.71 ;
      POLYGON 2.835 0.79 2.555 0.79 2.555 1.01 2.585 1.01 2.585 1.07 1.86 1.07 1.86 1.01 2.495 1.01 2.495 0.63 2.435 0.63 2.435 0.57 2.555 0.57 2.555 0.73 2.835 0.73 ;
      POLYGON 2.63 1.465 1.975 1.465 1.975 1.39 1.445 1.39 1.445 1.23 1.32 1.23 1.32 0.525 1.38 0.525 1.38 1.17 1.505 1.17 1.505 1.33 2.035 1.33 2.035 1.405 2.57 1.405 2.57 1.17 2.63 1.17 ;
      POLYGON 2.165 0.75 1.685 0.75 1.685 0.29 1.54 0.29 1.54 1.01 1.6 1.01 1.6 1.07 1.48 1.07 1.48 0.29 0.925 0.29 0.925 1.085 0.88 1.085 0.88 1.21 0.82 1.21 0.82 1.025 0.865 1.025 0.865 0.35 0.735 0.35 0.735 0.23 1.745 0.23 1.745 0.69 2.105 0.69 2.105 0.42 2.005 0.42 2.005 0.36 2.165 0.36 ;
      POLYGON 1.22 1.43 1.16 1.43 1.16 1.37 0.66 1.37 0.66 1.085 0.25 1.085 0.25 1.21 0.19 1.21 0.19 1.025 0.275 1.025 0.275 0.255 0.335 0.255 0.335 1.025 0.72 1.025 0.72 1.31 1.16 1.31 1.16 0.645 1.115 0.645 1.115 0.525 1.175 0.525 1.175 0.585 1.22 0.585 ;
  END
END TLATNTSCAX3

MACRO TLATNTSCAX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX4 0 0 ;
  SIZE 4.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.575 1.005 0.815 1.175 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.435 0.815 0.925 0.905 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.175 1.06 0.14 1.06 0.14 1.15 0.06 1.15 0.06 0.98 0.095 0.98 0.095 0.685 0.175 0.685 ;
    END
  END E
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.409 LAYER Metal1 ;
    ANTENNADIFFAREA 2.383225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.2565 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.39181275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 75.0643275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.915 1.385 3.855 1.385 3.855 0.73 3.55 0.73 3.55 1.03 3.505 1.03 3.505 1.385 3.445 1.385 3.445 0.97 3.49 0.97 3.49 0.73 3.46 0.73 3.46 0.585 3.445 0.585 3.445 0.465 3.52 0.465 3.52 0.6 3.54 0.6 3.54 0.67 3.855 0.67 3.855 0.465 3.915 0.465 ;
    END
  END ECK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 1.77 0 1.77 0 1.65 0.54 1.65 0.54 1.275 0.6 1.275 0.6 1.65 1.985 1.65 1.985 1.54 2.105 1.54 2.105 1.65 2.78 1.65 2.78 1.09 2.84 1.09 2.84 1.65 3.24 1.65 3.24 1.085 3.3 1.085 3.3 1.65 3.65 1.65 3.65 0.995 3.71 0.995 3.71 1.65 4.06 1.65 4.06 0.995 4.12 0.995 4.12 1.65 4.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.2 0.06 4.12 0.06 4.12 0.445 4.06 0.445 4.06 0.06 3.71 0.06 3.71 0.445 3.65 0.445 3.65 0.06 3.3 0.06 3.3 0.445 3.24 0.445 3.24 0.06 2.765 0.06 2.765 0.605 2.705 0.605 2.705 0.06 2.07 0.06 2.07 0.605 1.95 0.605 1.95 0.545 2.01 0.545 2.01 0.06 0.57 0.06 0.57 0.495 0.63 0.495 0.63 0.555 0.51 0.555 0.51 0.06 0.175 0.06 0.175 0.585 0.115 0.585 0.115 0.06 0 0.06 0 -0.06 4.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.39 0.87 3.255 0.87 3.255 0.985 3.095 0.985 3.095 1.385 3.035 1.385 3.035 0.925 3.195 0.925 3.195 0.605 3.015 0.605 3.015 0.485 3.075 0.485 3.075 0.545 3.255 0.545 3.255 0.81 3.39 0.81 ;
      POLYGON 3.095 0.825 3.035 0.825 3.035 0.765 2.545 0.765 2.545 0.41 2.245 0.41 2.245 0.705 2.28 0.705 2.28 1.025 2.34 1.025 2.34 1.085 2.22 1.085 2.22 0.765 1.765 0.765 1.765 0.375 1.445 0.375 1.445 1.175 1.385 1.175 1.385 0.315 1.825 0.315 1.825 0.705 2.185 0.705 2.185 0.35 2.605 0.35 2.605 0.705 3.095 0.705 ;
      POLYGON 2.935 0.925 2.585 0.925 2.585 1.245 1.945 1.245 1.945 1.19 1.885 1.19 1.885 1.13 2.005 1.13 2.005 1.185 2.525 1.185 2.525 0.925 2.385 0.925 2.385 0.51 2.445 0.51 2.445 0.865 2.935 0.865 ;
      POLYGON 2.68 1.405 1.545 1.405 1.545 0.57 1.665 0.57 1.665 0.63 1.605 0.63 1.605 1.285 1.65 1.285 1.65 1.345 2.68 1.345 ;
      POLYGON 2.12 0.945 1.825 0.945 1.825 1.03 1.705 1.03 1.705 0.95 1.745 0.95 1.745 0.865 2.12 0.865 ;
      POLYGON 1.445 1.395 1.385 1.395 1.385 1.335 1.225 1.335 1.225 0.39 0.925 0.39 0.925 0.715 0.335 0.715 0.335 1.31 0.2 1.31 0.2 1.25 0.275 1.25 0.275 0.655 0.32 0.655 0.32 0.49 0.38 0.49 0.38 0.655 0.865 0.655 0.865 0.33 1.285 0.33 1.285 1.275 1.445 1.275 ;
      POLYGON 1.125 1.06 1.085 1.06 1.085 1.335 0.805 1.335 0.805 1.395 0.745 1.395 0.745 1.275 1.025 1.275 1.025 0.49 1.085 0.49 1.085 0.94 1.125 0.94 ;
  END
END TLATNTSCAX4

MACRO TLATNTSCAX6
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX6 0 0 ;
  SIZE 5 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.7971 LAYER Metal1 ;
    ANTENNADIFFAREA 3.133475 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.380475 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.3516 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 58.02483725 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.74 0.66 4.695 0.66 4.695 0.76 4.74 0.76 4.74 1.37 4.68 1.37 4.68 0.82 4.33 0.82 4.33 1.37 4.27 1.37 4.27 0.82 3.94 0.82 3.94 0.92 3.92 0.92 3.92 1.37 3.86 1.37 3.86 0.35 3.92 0.35 3.92 0.76 4.27 0.76 4.27 0.35 4.33 0.35 4.33 0.76 4.635 0.76 4.635 0.6 4.68 0.6 4.68 0.35 4.74 0.35 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.66 0.45 0.74 0.95 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.46 0.45 0.54 0.95 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.2 0.895 0.035 0.895 0.035 0.815 0.08 0.815 0.08 0.48 0.2 0.48 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 1.77 0 1.77 0 1.65 0.525 1.65 0.525 1.21 0.585 1.21 0.585 1.65 2 1.65 2 1.49 2.12 1.49 2.12 1.55 2.06 1.55 2.06 1.65 2.835 1.65 2.835 1.01 2.895 1.01 2.895 1.65 3.245 1.65 3.245 1.25 3.305 1.25 3.305 1.65 3.655 1.65 3.655 1.25 3.715 1.25 3.715 1.65 4.065 1.65 4.065 0.92 4.125 0.92 4.125 1.65 4.475 1.65 4.475 0.92 4.535 0.92 4.535 1.65 5 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5 0.06 4.535 0.06 4.535 0.66 4.475 0.66 4.475 0.06 4.125 0.06 4.125 0.66 4.065 0.66 4.065 0.06 3.715 0.06 3.715 0.47 3.655 0.47 3.655 0.06 3.045 0.06 3.045 0.17 2.925 0.17 2.925 0.06 2.12 0.06 2.12 0.17 2 0.17 2 0.06 0.585 0.06 0.585 0.35 0.525 0.35 0.525 0.06 0.155 0.06 0.155 0.35 0.095 0.35 0.095 0.06 0 0.06 0 -0.06 5 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.76 1.1 3.51 1.1 3.51 1.37 3.45 1.37 3.45 1.1 3.1 1.1 3.1 1.37 3.04 1.37 3.04 1.04 3.7 1.04 3.7 0.74 3.495 0.74 3.495 0.56 3.295 0.56 3.295 0.44 3.355 0.44 3.355 0.5 3.555 0.5 3.555 0.68 3.76 0.68 ;
      POLYGON 3.6 0.9 3.44 0.9 3.44 0.94 2.975 0.94 2.975 0.75 2.515 0.75 2.515 1.01 2.575 1.01 2.575 1.07 2.455 1.07 2.455 0.88 1.99 0.88 1.99 0.82 2.455 0.82 2.455 0.69 2.69 0.69 2.69 0.53 2.81 0.53 2.81 0.59 2.75 0.59 2.75 0.69 3.035 0.69 3.035 0.88 3.38 0.88 3.38 0.84 3.6 0.84 ;
      POLYGON 3.28 0.78 3.22 0.78 3.22 0.72 3.135 0.72 3.135 0.59 2.91 0.59 2.91 0.43 2.44 0.43 2.44 0.525 2.325 0.525 2.325 0.72 1.89 0.72 1.89 1.01 2.355 1.01 2.355 1.07 1.83 1.07 1.83 0.72 1.77 0.72 1.77 0.66 2.265 0.66 2.265 0.465 2.38 0.465 2.38 0.37 2.97 0.37 2.97 0.53 3.195 0.53 3.195 0.66 3.28 0.66 ;
      POLYGON 2.86 0.91 2.735 0.91 2.735 1.23 1.605 1.23 1.605 1.1 1.45 1.1 1.45 0.56 1.39 0.56 1.39 0.5 1.51 0.5 1.51 1.04 1.665 1.04 1.665 1.17 2.675 1.17 2.675 0.85 2.86 0.85 ;
      POLYGON 2.28 0.365 1.67 0.365 1.67 0.82 1.73 0.82 1.73 0.94 1.67 0.94 1.67 0.88 1.61 0.88 1.61 0.365 1.385 0.365 1.385 0.315 0.905 0.315 0.905 1.145 0.965 1.145 0.965 1.205 0.845 1.205 0.845 0.255 1.445 0.255 1.445 0.305 2.28 0.305 ;
      POLYGON 1.35 1.365 0.685 1.365 0.685 1.11 0.305 1.11 0.305 1.205 0.185 1.205 0.185 1.145 0.245 1.145 0.245 1.05 0.3 1.05 0.3 0.255 0.36 0.255 0.36 1.05 0.745 1.05 0.745 1.305 1.23 1.305 1.23 1.045 1.215 1.045 1.215 0.47 1.275 0.47 1.275 0.985 1.29 0.985 1.29 1.075 1.35 1.075 ;
  END
END TLATNTSCAX6

MACRO TLATNTSCAX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNTSCAX8 0 0 ;
  SIZE 5.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN ECK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.928 LAYER Metal1 ;
    ANTENNADIFFAREA 3.307875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.438075 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.683787 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 53.2922445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.97 1.405 4.91 1.405 4.91 1.02 4.56 1.02 4.56 1.405 4.5 1.405 4.5 1.02 4.15 1.02 4.15 1.405 4.09 1.405 4.09 1.02 3.74 1.02 3.74 1.405 3.68 1.405 3.68 1.11 3.66 1.11 3.66 0.96 3.68 0.96 3.68 0.515 3.74 0.515 3.74 0.96 4.91 0.96 4.91 0.62 4.135 0.62 4.135 0.605 4.06 0.605 4.06 0.545 4.18 0.545 4.18 0.56 4.47 0.56 4.47 0.545 4.59 0.545 4.59 0.56 4.91 0.56 4.91 0.5 4.97 0.5 ;
    END
  END ECK
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.755 0.935 0.675 0.935 0.675 0.73 0.66 0.73 0.66 0.45 0.74 0.45 0.74 0.6 0.755 0.6 ;
    END
  END CK
  PIN SE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 0.73 0.525 0.73 0.525 0.935 0.445 0.935 0.445 0.45 0.54 0.45 ;
    END
  END SE
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.27777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.145 0.545 0.14 0.545 0.14 0.895 0.06 0.895 0.06 0.425 0.145 0.425 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.2 1.77 0 1.77 0 1.65 0.54 1.65 0.54 1.255 0.48 1.255 0.48 1.195 0.6 1.195 0.6 1.65 1.785 1.65 1.785 1.31 1.725 1.31 1.725 1.25 1.845 1.25 1.845 1.65 2.655 1.65 2.655 1.095 2.715 1.095 2.715 1.65 3.065 1.65 3.065 1.285 3.125 1.285 3.125 1.65 3.475 1.65 3.475 1.285 3.535 1.285 3.535 1.65 3.885 1.65 3.885 1.12 3.945 1.12 3.945 1.65 4.295 1.65 4.295 1.12 4.355 1.12 4.355 1.65 4.705 1.65 4.705 1.12 4.765 1.12 4.765 1.65 5.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.2 0.06 4.765 0.06 4.765 0.46 4.705 0.46 4.705 0.06 4.355 0.06 4.355 0.46 4.295 0.46 4.295 0.06 3.945 0.06 3.945 0.46 3.885 0.46 3.885 0.06 3.52 0.06 3.52 0.46 3.46 0.46 3.46 0.06 2.88 0.06 2.88 0.515 2.82 0.515 2.82 0.06 2.02 0.06 2.02 0.35 1.9 0.35 1.9 0.29 1.96 0.29 1.96 0.06 0.57 0.06 0.57 0.35 0.51 0.35 0.51 0.06 0.14 0.06 0.14 0.35 0.08 0.35 0.08 0.06 0 0.06 0 -0.06 5.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.56 1.1 3.33 1.1 3.33 1.405 3.27 1.405 3.27 1.1 2.92 1.1 2.92 1.405 2.86 1.405 2.86 1.04 3.5 1.04 3.5 0.72 3.3 0.72 3.3 0.515 3.15 0.515 3.15 0.395 3.21 0.395 3.21 0.455 3.36 0.455 3.36 0.66 3.56 0.66 ;
      POLYGON 3.38 0.94 2.785 0.94 2.785 0.835 2.395 0.835 2.395 1.215 2.335 1.215 2.335 0.83 1.815 0.83 1.815 0.77 2.5 0.77 2.5 0.48 2.56 0.48 2.56 0.775 2.845 0.775 2.845 0.88 3.32 0.88 3.32 0.82 3.38 0.82 ;
      POLYGON 3.135 0.77 3.075 0.77 3.075 0.675 2.66 0.675 2.66 0.38 2.4 0.38 2.4 0.595 2.34 0.595 2.34 0.67 1.715 0.67 1.715 0.93 2.165 0.93 2.165 1.155 2.225 1.155 2.225 1.215 2.105 1.215 2.105 0.99 1.655 0.99 1.655 0.61 2.28 0.61 2.28 0.535 2.34 0.535 2.34 0.32 2.72 0.32 2.72 0.615 3.135 0.615 ;
      POLYGON 2.555 1.375 1.945 1.375 1.945 1.15 1.505 1.15 1.505 1.245 1.445 1.245 1.445 1.15 1.335 1.15 1.335 0.63 1.275 0.63 1.275 0.57 1.395 0.57 1.395 1.09 2.005 1.09 2.005 1.315 2.495 1.315 2.495 0.935 2.555 0.935 ;
      POLYGON 2.24 0.435 2.18 0.435 2.18 0.51 1.555 0.51 1.555 0.99 1.495 0.99 1.495 0.315 0.92 0.315 0.92 1.1 0.98 1.1 0.98 1.16 0.86 1.16 0.86 0.375 0.815 0.375 0.815 0.255 1.555 0.255 1.555 0.45 2.12 0.45 2.12 0.375 2.24 0.375 ;
      POLYGON 1.235 1.34 1.175 1.34 1.175 1.32 0.7 1.32 0.7 1.095 0.26 1.095 0.26 1.19 0.2 1.19 0.2 1.035 0.285 1.035 0.285 0.255 0.345 0.255 0.345 1.035 0.76 1.035 0.76 1.26 1.1 1.26 1.1 0.54 1.16 0.54 1.16 1.22 1.235 1.22 ;
  END
END TLATNTSCAX8

MACRO TLATNX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNX1 0 0 ;
  SIZE 3.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.788425 LAYER Metal1 ;
    ANTENNADIFFAREA 1.877125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.16875 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.598074 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 81.7244445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.175 1.29 3.095 1.29 3.095 0.515 3.035 0.515 3.035 0.435 3.07 0.435 3.07 0.395 3.175 0.395 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.788425 LAYER Metal1 ;
    ANTENNADIFFAREA 1.877125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.16875 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.598074 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 81.7244445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.46 0.54 2.54 1.34 ;
    END
  END QN
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.165 1.085 2.115 1.085 2.115 1.23 2.035 1.23 2.035 0.78 2.115 0.78 2.115 1.005 2.165 1.005 ;
    END
  END GN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.53 0.98 0.26 0.98 0.26 0.785 0.34 0.785 0.34 0.9 0.45 0.9 0.45 0.785 0.53 0.785 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 1.77 0 1.77 0 1.65 0.46 1.65 0.46 1.24 0.52 1.24 0.52 1.65 1.29 1.65 1.29 1.51 1.35 1.51 1.35 1.65 2.255 1.65 2.255 1.185 2.315 1.185 2.315 1.65 2.865 1.65 2.865 0.9 2.925 0.9 2.925 1.65 3.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.4 0.06 2.925 0.06 2.925 0.515 2.865 0.515 2.865 0.06 2.295 0.06 2.295 0.52 2.235 0.52 2.235 0.06 1.295 0.06 1.295 0.525 1.235 0.525 1.235 0.06 0.49 0.06 0.49 0.525 0.43 0.525 0.43 0.06 0 0.06 0 -0.06 3.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.995 0.785 2.72 0.785 2.72 1.29 2.66 1.29 2.66 0.535 2.72 0.535 2.72 0.725 2.995 0.725 ;
      POLYGON 2.36 0.82 2.3 0.82 2.3 0.68 2.075 0.68 2.075 0.44 1.585 0.44 1.585 1.165 1.525 1.165 1.525 0.945 1.255 0.945 1.255 1.005 1.195 1.005 1.195 0.885 1.525 0.885 1.525 0.525 1.44 0.525 1.44 0.38 2.135 0.38 2.135 0.62 2.36 0.62 ;
      POLYGON 1.935 1.385 0.79 1.385 0.79 0.945 0.875 0.945 0.875 0.685 0.335 0.685 0.335 0.625 0.935 0.625 0.935 1.005 0.85 1.005 0.85 1.325 1.875 1.325 1.875 0.54 1.935 0.54 ;
      POLYGON 1.425 0.785 1.095 0.785 1.095 1.165 1.01 1.165 1.01 1.225 0.95 1.225 0.95 1.105 1.035 1.105 1.035 0.525 0.74 0.525 0.74 0.405 0.8 0.405 0.8 0.465 1.095 0.465 1.095 0.725 1.365 0.725 1.365 0.665 1.425 0.665 ;
      POLYGON 0.775 0.845 0.69 0.845 0.69 1.14 0.285 1.14 0.285 1.2 0.225 1.2 0.225 1.14 0.1 1.14 0.1 0.465 0.225 0.465 0.225 0.405 0.285 0.405 0.285 0.525 0.16 0.525 0.16 1.08 0.63 1.08 0.63 0.785 0.775 0.785 ;
  END
END TLATNX1

MACRO TLATNX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNX2 0 0 ;
  SIZE 3.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 0.06 3.37 0.06 3.37 0.44 3.31 0.44 3.31 0.06 2.935 0.06 2.935 0.44 2.875 0.44 2.875 0.06 2.525 0.06 2.525 0.44 2.465 0.44 2.465 0.06 2.115 0.06 2.115 0.17 1.995 0.17 1.995 0.06 1.335 0.06 1.335 0.425 1.275 0.425 1.275 0.06 0.465 0.06 0.465 0.425 0.405 0.425 0.405 0.06 0 0.06 0 -0.06 3.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 1.77 0 1.77 0 1.65 0.41 1.65 0.41 1.155 0.47 1.155 0.47 1.65 1.275 1.65 1.275 1.54 1.395 1.54 1.395 1.65 1.995 1.65 1.995 0.995 2.055 0.995 2.055 1.65 2.465 1.65 2.465 0.9 2.525 0.9 2.525 1.65 2.875 1.65 2.875 0.9 2.935 0.9 2.935 1.65 3.31 1.65 3.31 0.9 3.37 0.9 3.37 1.65 3.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.565 0.765 0.515 0.765 0.515 0.895 0.195 0.895 0.195 0.815 0.435 0.815 0.435 0.685 0.565 0.685 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.77777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.825 0.625 1.975 0.895 ;
    END
  END GN
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0246 LAYER Metal1 ;
    ANTENNADIFFAREA 2.1862 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.263475 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.6842205 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 59.53885575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.46 2.34 1.29 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.0246 LAYER Metal1 ;
    ANTENNADIFFAREA 2.1862 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.263475 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.6842205 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 59.53885575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.365 0.705 3.185 0.705 3.185 1.29 3.105 1.29 3.105 0.46 3.185 0.46 3.185 0.625 3.365 0.625 ;
    END
  END Q
  OBS
    LAYER Metal1 ;
      POLYGON 3.005 0.71 2.73 0.71 2.73 1.29 2.67 1.29 2.67 0.46 2.73 0.46 2.73 0.65 3.005 0.65 ;
      POLYGON 2.16 0.74 2.1 0.74 2.1 0.365 1.565 0.365 1.565 1.155 1.63 1.155 1.63 1.215 1.505 1.215 1.505 0.95 1.31 0.95 1.31 1.01 1.25 1.01 1.25 0.89 1.505 0.89 1.505 0.305 2.16 0.305 ;
      POLYGON 1.88 0.525 1.725 0.525 1.725 0.995 1.85 0.995 1.85 1.405 0.775 1.405 0.775 1.025 0.93 1.025 0.93 0.645 0.665 0.645 0.665 0.585 0.335 0.585 0.335 0.645 0.275 0.645 0.275 0.525 0.99 0.525 0.99 1.085 0.835 1.085 0.835 1.345 1.79 1.345 1.79 1.055 1.665 1.055 1.665 0.465 1.88 0.465 ;
      POLYGON 1.405 0.64 1.15 0.64 1.15 1.245 0.935 1.245 0.935 1.185 1.09 1.185 1.09 0.425 0.72 0.425 0.72 0.305 0.78 0.305 0.78 0.365 1.15 0.365 1.15 0.58 1.405 0.58 ;
      POLYGON 0.83 0.925 0.675 0.925 0.675 1.055 0.265 1.055 0.265 1.18 0.205 1.18 0.205 1.055 0.035 1.055 0.035 0.365 0.2 0.365 0.2 0.305 0.26 0.305 0.26 0.425 0.095 0.425 0.095 0.995 0.615 0.995 0.615 0.865 0.83 0.865 ;
  END
END TLATNX2

MACRO TLATNX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNX4 0 0 ;
  SIZE 5.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8006 LAYER Metal1 ;
    ANTENNADIFFAREA 3.6152 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.46215 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.05993725 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 46.3550795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.18 0.575 2.925 0.575 2.925 1.005 3 1.005 3 1.34 2.94 1.34 2.94 1.065 2.765 1.065 2.765 1.085 2.59 1.085 2.59 1.34 2.53 1.34 2.53 1.005 2.865 1.005 2.865 0.575 2.65 0.575 2.65 0.455 2.71 0.455 2.71 0.515 3.12 0.515 3.12 0.455 3.18 0.455 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.8006 LAYER Metal1 ;
    ANTENNADIFFAREA 3.6152 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.46215 LAYER Metal1 ;
      ANTENNAMAXAREACAR 6.05993725 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 46.3550795 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.33 1.34 1.27 1.34 1.27 1.01 0.92 1.01 0.92 1.34 0.86 1.34 0.86 0.79 0.88 0.79 0.88 0.575 0.77 0.575 0.77 0.455 0.83 0.455 0.83 0.515 1.24 0.515 1.24 0.455 1.3 0.455 1.3 0.575 0.94 0.575 0.94 0.95 1.33 0.95 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.66 0.62 4.74 1.12 ;
    END
  END D
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.67 0.705 0.585 0.705 0.585 0.85 0.375 0.85 0.375 0.77 0.435 0.77 0.435 0.565 0.67 0.565 ;
    END
  END GN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.2 1.77 0 1.77 0 1.65 0.655 1.65 0.655 0.95 0.715 0.95 0.715 1.65 1.065 1.65 1.065 1.11 1.125 1.11 1.125 1.65 1.475 1.65 1.475 0.95 1.535 0.95 1.535 1.65 1.915 1.65 1.915 1.11 1.975 1.11 1.975 1.65 2.325 1.65 2.325 0.95 2.385 0.95 2.385 1.65 2.735 1.65 2.735 1.22 2.795 1.22 2.795 1.65 3.195 1.65 3.195 0.95 3.255 0.95 3.255 1.65 3.605 1.65 3.605 1.25 3.725 1.25 3.725 1.31 3.665 1.31 3.665 1.65 4.66 1.65 4.66 1.22 4.72 1.22 4.72 1.65 5.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.2 0.06 4.69 0.06 4.69 0.2 4.63 0.2 4.63 0.06 3.97 0.06 3.97 0.2 3.91 0.2 3.91 0.06 3.445 0.06 3.445 0.17 3.325 0.17 3.325 0.06 2.975 0.06 2.975 0.17 2.855 0.17 2.855 0.06 2.505 0.06 2.505 0.17 2.385 0.17 2.385 0.06 2.035 0.06 2.035 0.17 1.915 0.17 1.915 0.06 1.565 0.06 1.565 0.17 1.445 0.17 1.445 0.06 1.095 0.06 1.095 0.17 0.975 0.17 0.975 0.06 0.51 0.06 0.51 0.2 0.45 0.2 0.45 0.06 0 0.06 0 -0.06 5.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.985 0.52 4.925 0.52 4.925 1.245 4.865 1.245 4.865 0.52 4.56 0.52 4.56 0.84 4.44 0.84 4.44 0.46 4.985 0.46 ;
      POLYGON 4.91 0.35 4.85 0.35 4.85 0.36 4.12 0.36 4.12 0.885 4.18 0.885 4.18 0.945 4.06 0.945 4.06 0.36 3.75 0.36 3.75 0.355 0.67 0.355 0.67 0.36 0.275 0.36 0.275 0.95 0.48 0.95 0.48 1.07 0.42 1.07 0.42 1.01 0.215 1.01 0.215 0.3 0.61 0.3 0.61 0.295 3.81 0.295 3.81 0.3 4.27 0.3 4.27 0.16 4.39 0.16 4.39 0.3 4.79 0.3 4.79 0.29 4.91 0.29 ;
      POLYGON 4.34 1.245 4.28 1.245 4.28 1.105 3.825 1.105 3.825 0.98 3.59 0.98 3.59 0.86 3.65 0.86 3.65 0.92 3.885 0.92 3.885 1.045 4.28 1.045 4.28 0.545 4.22 0.545 4.22 0.485 4.34 0.485 ;
      POLYGON 3.96 0.76 3.9 0.76 3.9 0.7 3.49 0.7 3.49 1.34 3.43 1.34 3.43 0.735 3.025 0.735 3.025 0.675 3.43 0.675 3.43 0.64 3.59 0.64 3.59 0.455 3.65 0.455 3.65 0.64 3.96 0.64 ;
      POLYGON 2.24 0.575 1.77 0.575 1.77 0.95 2.18 0.95 2.18 1.34 2.12 1.34 2.12 1.01 1.77 1.01 1.77 1.34 1.71 1.34 1.71 0.85 1.275 0.85 1.275 0.79 1.71 0.79 1.71 0.455 1.77 0.455 1.77 0.515 2.18 0.515 2.18 0.455 2.24 0.455 ;
  END
END TLATNX4

MACRO TLATNXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATNXL 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.72005 LAYER Metal1 ;
    ANTENNADIFFAREA 1.6228 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1296 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.27199075 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 103.3680555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.06 0.405 3.14 1.02 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.76925 LAYER Metal1 ;
    ANTENNADIFFAREA 1.6228 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1296 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.65162025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 104.97685175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.355 1.385 2.26 1.385 2.26 0.405 2.34 0.405 2.34 1.265 2.355 1.265 ;
    END
  END QN
  PIN GN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.06 0.76 2.14 1.26 ;
    END
  END GN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.48 1.11 0.34 1.11 0.34 1.12 0.26 1.12 0.26 0.955 0.4 0.955 0.4 0.76 0.48 0.76 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 1.77 0 1.77 0 1.65 0.345 1.65 0.345 1.51 0.405 1.51 0.405 1.65 1.3 1.65 1.3 1.51 1.36 1.51 1.36 1.65 2.09 1.65 2.09 1.36 2.15 1.36 2.15 1.65 2.83 1.65 2.83 0.995 2.89 0.995 2.89 1.65 3.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 0.06 2.89 0.06 2.89 0.5 2.83 0.5 2.83 0.06 2 0.06 2 0.5 1.94 0.5 1.94 0.06 1.23 0.06 1.23 0.495 1.17 0.495 1.17 0.06 0.375 0.06 0.375 0.495 0.315 0.495 0.315 0.06 0 0.06 0 -0.06 3.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.96 0.68 2.705 0.68 2.705 1.02 2.625 1.02 2.625 0.405 2.705 0.405 2.705 0.6 2.96 0.6 ;
      POLYGON 2.22 0.3 2.16 0.3 2.16 0.66 1.78 0.66 1.78 0.305 1.52 0.305 1.52 1.125 1.595 1.125 1.595 1.245 1.535 1.245 1.535 1.185 1.46 1.185 1.46 0.875 1.34 0.875 1.34 0.935 1.28 0.935 1.28 0.815 1.46 0.815 1.46 0.495 1.375 0.495 1.375 0.245 1.84 0.245 1.84 0.6 2.1 0.6 2.1 0.24 2.22 0.24 ;
      POLYGON 1.94 1.48 1.88 1.48 1.88 1.42 1.715 1.42 1.715 1.41 0.8 1.41 0.8 0.66 0.3 0.66 0.3 0.715 0.24 0.715 0.24 0.595 0.3 0.595 0.3 0.6 0.86 0.6 0.86 0.97 0.96 0.97 0.96 0.91 1.02 0.91 1.02 1.03 0.86 1.03 0.86 1.35 1.695 1.35 1.695 1.025 1.62 1.025 1.62 0.405 1.68 0.405 1.68 0.965 1.755 0.965 1.755 1.36 1.94 1.36 ;
      POLYGON 1.36 0.715 1.18 0.715 1.18 1.19 1.02 1.19 1.02 1.25 0.96 1.25 0.96 1.13 1.12 1.13 1.12 0.715 1.01 0.715 1.01 0.5 0.65 0.5 0.65 0.38 0.71 0.38 0.71 0.44 1.07 0.44 1.07 0.655 1.3 0.655 1.3 0.595 1.36 0.595 ;
      POLYGON 0.7 1.055 0.64 1.055 0.64 1.28 0.17 1.28 0.17 1.34 0.08 1.34 0.08 0.4 0.14 0.4 0.14 1.22 0.58 1.22 0.58 0.995 0.7 0.995 ;
  END
END TLATNXL

MACRO TLATSRX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATSRX1 0 0 ;
  SIZE 3.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.97815 LAYER Metal1 ;
    ANTENNADIFFAREA 2.189575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.16875 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.72237025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 89.92 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.94 1.07 0.88 1.07 0.88 0.73 0.86 0.73 0.86 0.6 0.88 0.6 0.88 0.41 0.94 0.41 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.02035 LAYER Metal1 ;
    ANTENNADIFFAREA 2.189575 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.16875 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.9724445 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 91.2355555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.305 1.29 0.225 1.29 0.225 0.54 0.06 0.54 0.06 0.41 0.305 0.41 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.47 1.155 3.26 1.155 3.26 0.845 3.39 0.845 3.39 0.785 3.47 0.785 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.43 0.96 2.025 0.96 2.025 0.785 2.105 0.785 2.105 0.815 2.43 0.815 ;
    END
  END RN
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.765 0.895 1.68 0.895 1.68 1.23 1.6 1.23 1.6 0.815 1.765 0.815 ;
    END
  END G
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.34 1.09 1.26 1.09 1.26 0.92 1.2 0.92 1.2 0.84 1.26 0.84 1.26 0.65 1.34 0.65 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 1.77 0 1.77 0 1.65 0.475 1.65 0.475 0.9 0.535 0.9 0.535 1.65 1.085 1.65 1.085 1.19 1.145 1.19 1.145 1.65 1.54 1.65 1.54 1.51 1.6 1.51 1.6 1.65 2.12 1.65 2.12 1.51 2.18 1.51 2.18 1.65 2.52 1.65 2.52 1.4 2.58 1.4 2.58 1.65 3.405 1.65 3.405 1.54 3.525 1.54 3.525 1.65 3.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.8 0.06 3.525 0.06 3.525 0.525 3.465 0.525 3.465 0.06 2.46 0.06 2.46 0.365 2.34 0.365 2.34 0.305 2.4 0.305 2.4 0.06 1.145 0.06 1.145 0.39 1.085 0.39 1.085 0.06 0.535 0.06 0.535 0.52 0.475 0.52 0.475 0.06 0 0.06 0 -0.06 3.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.745 1.36 3.225 1.36 3.225 1.445 3.105 1.445 3.105 1.36 2.91 1.36 2.91 0.685 1.925 0.685 1.925 1.215 1.865 1.215 1.865 0.46 1.985 0.46 1.985 0.52 1.925 0.52 1.925 0.625 2.97 0.625 2.97 1.3 3.745 1.3 ;
      POLYGON 3.73 1.135 3.67 1.135 3.67 0.685 3.29 0.685 3.29 0.745 3.23 0.745 3.23 0.625 3.67 0.625 3.67 0.43 3.73 0.43 ;
      POLYGON 3.13 1.135 3.07 1.135 3.07 0.525 2.18 0.525 2.18 0.31 1.37 0.31 1.37 0.25 2.24 0.25 2.24 0.465 3.07 0.465 3.07 0.405 3.13 0.405 ;
      POLYGON 2.81 1.125 2.77 1.125 2.77 1.3 2.255 1.3 2.255 1.22 2.69 1.22 2.69 1.045 2.81 1.045 ;
      POLYGON 2.59 1.12 2.155 1.12 2.155 1.41 1.305 1.41 1.305 1.19 1.44 1.19 1.44 0.55 1.1 0.55 1.1 0.7 1.04 0.7 1.04 0.49 1.465 0.49 1.465 0.41 1.525 0.41 1.525 0.55 1.5 0.55 1.5 1.25 1.365 1.25 1.365 1.35 2.095 1.35 2.095 1.06 2.53 1.06 2.53 0.91 2.59 0.91 ;
      POLYGON 0.74 1.02 0.66 1.02 0.66 0.8 0.405 0.8 0.405 0.72 0.66 0.72 0.66 0.54 0.74 0.54 ;
  END
END TLATSRX1

MACRO TLATSRX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATSRX2 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.574 LAYER Metal1 ;
    ANTENNADIFFAREA 2.894825 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.263475 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.76942775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 76.2766865 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.54 0.92 4.38 0.92 4.38 0.935 4.335 0.935 4.335 1.345 4.275 1.345 4.275 0.875 4.32 0.875 4.32 0.62 4.275 0.62 4.275 0.5 4.335 0.5 4.335 0.56 4.38 0.56 4.38 0.79 4.54 0.79 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.574 LAYER Metal1 ;
    ANTENNADIFFAREA 2.894825 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.263475 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.76942775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 76.2766865 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.765 0.705 3.635 0.705 3.635 0.685 3.535 0.685 3.535 0.91 3.515 0.91 3.515 1.345 3.455 1.345 3.455 0.85 3.475 0.85 3.475 0.535 3.455 0.535 3.455 0.415 3.515 0.415 3.515 0.475 3.535 0.475 3.535 0.625 3.765 0.625 ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.285 1.085 3.115 1.085 3.115 1.125 3.035 1.125 3.035 0.795 3.155 0.795 3.155 1.005 3.285 1.005 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 1.11 1.86 1.11 1.86 0.985 1.565 0.985 1.565 0.905 1.94 0.905 ;
    END
  END RN
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.7 1 0.62 1 0.62 0.92 0.46 0.92 0.46 0.66 0.7 0.66 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 2.26 0.53 2.34 1.03 ;
    END
  END G
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.46 1.65 0.46 1.26 0.52 1.26 0.52 1.65 1.475 1.65 1.475 1.54 1.595 1.54 1.595 1.65 1.905 1.65 1.905 1.51 1.965 1.51 1.965 1.65 2.62 1.65 2.62 1.51 2.68 1.51 2.68 1.65 3.16 1.65 3.16 1.225 3.22 1.225 3.22 1.65 3.66 1.65 3.66 0.955 3.72 0.955 3.72 1.65 4.07 1.65 4.07 0.955 4.13 0.955 4.13 1.65 4.48 1.65 4.48 1.02 4.54 1.02 4.54 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 4.54 0.06 4.54 0.48 4.48 0.48 4.48 0.06 4.13 0.06 4.13 0.48 4.07 0.48 4.07 0.06 3.72 0.06 3.72 0.48 3.66 0.48 3.66 0.06 3.22 0.06 3.22 0.535 3.16 0.535 3.16 0.06 1.895 0.06 1.895 0.25 1.775 0.25 1.775 0.19 1.835 0.19 1.835 0.06 0.405 0.06 0.405 0.34 0.465 0.34 0.465 0.4 0.345 0.4 0.345 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.22 0.775 3.925 0.775 3.925 1.345 3.865 1.345 3.865 0.5 3.925 0.5 3.925 0.715 4.22 0.715 ;
      POLYGON 3.375 0.75 3.255 0.75 3.255 0.695 2.935 0.695 2.935 1.345 2.875 1.345 2.875 0.695 2.85 0.695 2.85 0.22 2.055 0.22 2.055 0.41 1.615 0.41 1.615 0.24 1.5 0.24 1.5 0.18 1.675 0.18 1.675 0.35 1.995 0.35 1.995 0.16 2.91 0.16 2.91 0.635 3.375 0.635 ;
      POLYGON 2.775 1.41 1.075 1.41 1.075 1.005 1.09 1.005 1.09 0.965 1.18 0.965 1.18 0.335 1.24 0.335 1.24 1.025 1.15 1.025 1.15 1.065 1.135 1.065 1.135 1.35 2.715 1.35 2.715 0.875 2.775 0.875 ;
      POLYGON 2.5 1.19 2.13 1.19 2.13 1.25 2.07 1.25 2.07 1.19 2.04 1.19 2.04 0.725 1.34 0.725 1.34 0.235 1.08 0.235 1.08 0.865 1.02 0.865 1.02 0.56 0.36 0.56 0.36 0.625 0.3 0.625 0.3 0.5 1.02 0.5 1.02 0.175 1.4 0.175 1.4 0.665 2.1 0.665 2.1 1.13 2.44 1.13 2.44 0.43 2.335 0.43 2.335 0.31 2.395 0.31 2.395 0.37 2.5 0.37 ;
      RECT 1.25 1.125 1.76 1.205 ;
      POLYGON 0.92 0.73 0.86 0.73 0.86 1.16 0.285 1.16 0.285 1.22 0.225 1.22 0.225 1.16 0.14 1.16 0.14 0.335 0.2 0.335 0.2 1.1 0.8 1.1 0.8 0.67 0.92 0.67 ;
  END
END TLATSRX2

MACRO TLATSRX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATSRX4 0 0 ;
  SIZE 7.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6698 LAYER Metal1 ;
    ANTENNADIFFAREA 5.219875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.46215 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.940712 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 59.363843 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.42 0.735 4.16 0.735 4.16 0.995 4.22 0.995 4.22 1.055 3.6 1.055 3.6 0.995 3.66 0.995 3.66 0.465 3.72 0.465 3.72 0.79 3.74 0.79 3.74 0.995 4.1 0.995 4.1 0.675 4.36 0.675 4.36 0.465 4.42 0.465 ;
    END
  END QN
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04635 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.33980575 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 4.775 0.815 5.52 0.895 ;
    END
  END SN
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 78.287037 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 5.835 0.37 5.775 0.37 5.775 0.41 5.335 0.41 5.335 0.365 4.96 0.365 4.96 0.555 4.52 0.555 4.52 0.365 4.26 0.365 4.26 0.575 3.82 0.575 3.82 0.365 3.56 0.365 3.56 0.605 3.18 0.605 3.18 0.365 2.92 0.365 2.92 0.605 2.54 0.605 2.54 0.365 2.28 0.365 2.28 0.605 1.9 0.605 1.9 0.365 1.64 0.365 1.64 0.605 1.26 0.605 1.26 0.365 1 0.365 1 0.66 0.74 0.66 0.74 0.73 0.735 0.73 0.735 0.78 0.66 0.78 0.66 0.6 0.94 0.6 0.94 0.305 1.32 0.305 1.32 0.545 1.58 0.545 1.58 0.305 1.96 0.305 1.96 0.545 2.22 0.545 2.22 0.305 2.6 0.305 2.6 0.545 2.86 0.545 2.86 0.305 3.24 0.305 3.24 0.545 3.5 0.545 3.5 0.305 3.88 0.305 3.88 0.515 4.2 0.515 4.2 0.305 4.58 0.305 4.58 0.495 4.9 0.495 4.9 0.305 5.395 0.305 5.395 0.35 5.715 0.35 5.715 0.31 5.835 0.31 ;
    END
  END RN
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.4 0.895 0.03 0.895 0.03 0.795 0.28 0.795 0.28 0.685 0.4 0.685 ;
    END
  END G
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.14 0.92 7.06 0.92 7.06 0.91 6.82 0.91 6.82 0.66 6.9 0.66 6.9 0.79 7.14 0.79 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.6698 LAYER Metal1 ;
    ANTENNADIFFAREA 5.219875 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.46215 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.940712 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 59.363843 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.055 1.07 1.055 1.07 0.995 1.1 0.995 1.1 0.465 1.16 0.465 1.16 0.79 1.34 0.79 1.34 0.995 1.74 0.995 1.74 0.465 1.8 0.465 ;
    END
  END Q
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.6 1.77 0 1.77 0 1.65 0.295 1.65 0.295 1.06 0.355 1.06 0.355 1.65 0.865 1.65 0.865 1.51 0.925 1.51 0.925 1.65 1.305 1.65 1.305 1.315 1.425 1.315 1.425 1.375 1.365 1.375 1.365 1.65 1.995 1.65 1.995 1.315 2.115 1.315 2.115 1.375 2.055 1.375 2.055 1.65 2.585 1.65 2.585 1.315 2.705 1.315 2.705 1.375 2.645 1.375 2.645 1.65 3.225 1.65 3.225 1.315 3.345 1.315 3.345 1.375 3.285 1.375 3.285 1.65 3.865 1.65 3.865 1.315 3.985 1.315 3.985 1.375 3.925 1.375 3.925 1.65 4.49 1.65 4.49 1.315 4.61 1.315 4.61 1.375 4.55 1.375 4.55 1.65 5.09 1.65 5.09 1.51 5.15 1.51 5.15 1.65 5.525 1.65 5.525 1.51 5.585 1.51 5.585 1.65 5.92 1.65 5.92 1.54 6.04 1.54 6.04 1.65 6.895 1.65 6.895 1.18 6.955 1.18 6.955 1.65 7.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 7.6 0.06 6.955 0.06 6.955 0.34 7.015 0.34 7.015 0.4 6.895 0.4 6.895 0.06 5.615 0.06 5.615 0.25 5.495 0.25 5.495 0.19 5.555 0.19 5.555 0.06 4.8 0.06 4.8 0.395 4.68 0.395 4.68 0.335 4.74 0.335 4.74 0.06 4.1 0.06 4.1 0.415 3.98 0.415 3.98 0.355 4.04 0.355 4.04 0.06 3.4 0.06 3.4 0.445 3.34 0.445 3.34 0.06 2.76 0.06 2.76 0.445 2.7 0.445 2.7 0.06 2.12 0.06 2.12 0.445 2.06 0.445 2.06 0.06 1.48 0.06 1.48 0.445 1.42 0.445 1.42 0.06 0.84 0.06 0.84 0.445 0.78 0.445 0.78 0.06 0 0.06 0 -0.06 7.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 7.46 1.205 7.4 1.205 7.4 0.56 6.735 0.56 6.735 0.555 6.465 0.555 6.465 0.37 6.405 0.37 6.405 0.31 6.525 0.31 6.525 0.495 6.795 0.495 6.795 0.5 7.315 0.5 7.315 0.44 7.375 0.44 7.375 0.5 7.46 0.5 ;
      POLYGON 7.3 1.08 6.72 1.08 6.72 1.395 5.13 1.395 5.13 1.215 0.5 1.215 0.5 0.585 0.44 0.585 0.44 0.465 0.5 0.465 0.5 0.525 0.56 0.525 0.56 1.155 5.19 1.155 5.19 1.335 6.34 1.335 6.34 1.055 6.215 1.055 6.215 0.815 6.275 0.815 6.275 0.995 6.4 0.995 6.4 1.335 6.66 1.335 6.66 0.735 6.6 0.735 6.6 0.675 6.72 0.675 6.72 1.02 7.24 1.02 7.24 0.915 7.3 0.915 ;
      POLYGON 6.56 1.205 6.5 1.205 6.5 0.895 6.375 0.895 6.375 0.715 5.22 0.715 5.22 0.655 6.29 0.655 6.29 0.465 6.35 0.465 6.35 0.655 6.435 0.655 6.435 0.835 6.56 0.835 ;
      RECT 5.685 1.155 6.24 1.235 ;
      POLYGON 5.88 0.95 5.68 0.95 5.68 1.055 5.35 1.055 5.35 1.115 5.29 1.115 5.29 1.055 4.615 1.055 4.615 0.895 4.395 0.895 4.395 0.835 4.615 0.835 4.615 0.655 5.06 0.655 5.06 0.465 5.12 0.465 5.12 0.715 4.675 0.715 4.675 0.995 5.62 0.995 5.62 0.89 5.88 0.89 ;
      POLYGON 3.08 1.055 2.96 1.055 2.96 0.995 3.02 0.995 3.02 0.765 2.47 0.765 2.47 1.055 2.35 1.055 2.35 0.995 2.41 0.995 2.41 0.765 1.9 0.765 1.9 0.705 2.38 0.705 2.38 0.465 2.44 0.465 2.44 0.705 3.02 0.705 3.02 0.465 3.08 0.465 ;
  END
END TLATSRX4

MACRO TLATSRXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATSRXL 0 0 ;
  SIZE 4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.034 LAYER Metal1 ;
    ANTENNADIFFAREA 2.161225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1296 LAYER Metal1 ;
      ANTENNAMAXAREACAR 15.6944445 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 117.22222225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.005 1.22 0.925 1.22 0.925 0.73 0.86 0.73 0.86 0.6 0.925 0.6 0.925 0.49 1.005 0.49 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.034 LAYER Metal1 ;
    ANTENNADIFFAREA 2.161225 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1296 LAYER Metal1 ;
      ANTENNAMAXAREACAR 15.6944445 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 117.22222225 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.325 1.02 0.245 1.02 0.245 0.73 0.06 0.73 0.06 0.6 0.245 0.6 0.245 0.54 0.325 0.54 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.67 1.06 3.54 1.06 3.54 1.185 3.46 1.185 3.46 0.98 3.59 0.98 3.59 0.815 3.67 0.815 ;
    END
  END D
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.37037025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.63 0.965 2.435 0.965 2.435 0.895 2.2 0.895 2.2 0.815 2.63 0.815 ;
    END
  END RN
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.61 1.94 1.11 ;
    END
  END G
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.06 1.265 1.06 1.265 0.96 1.435 0.96 1.435 0.815 1.6 0.815 ;
    END
  END SN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 1.77 0 1.77 0 1.65 0.525 1.65 0.525 1.285 0.585 1.285 0.585 1.65 1.21 1.65 1.21 1.51 1.27 1.51 1.27 1.65 1.73 1.65 1.73 1.51 1.79 1.51 1.79 1.65 2.39 1.65 2.39 1.51 2.45 1.51 2.45 1.65 2.79 1.65 2.79 1.405 2.85 1.405 2.85 1.65 3.605 1.65 3.605 1.54 3.725 1.54 3.725 1.65 4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4 0.06 3.725 0.06 3.725 0.555 3.665 0.555 3.665 0.06 2.675 0.06 2.675 0.395 2.555 0.395 2.555 0.335 2.615 0.335 2.615 0.06 1.21 0.06 1.21 0.495 1.27 0.495 1.27 0.555 1.15 0.555 1.15 0.06 0.555 0.06 0.555 0.635 0.495 0.635 0.495 0.06 0 0.06 0 -0.06 4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 3.945 1.365 3.425 1.365 3.425 1.475 3.305 1.475 3.305 1.365 3.11 1.365 3.11 0.715 2.1 0.715 2.1 1.22 2.04 1.22 2.04 0.49 2.16 0.49 2.16 0.55 2.1 0.55 2.1 0.655 3.17 0.655 3.17 1.305 3.945 1.305 ;
      POLYGON 3.93 1.14 3.87 1.14 3.87 0.715 3.49 0.715 3.49 0.75 3.43 0.75 3.43 0.63 3.49 0.63 3.49 0.655 3.87 0.655 3.87 0.46 3.93 0.46 ;
      POLYGON 3.33 1.14 3.27 1.14 3.27 0.555 2.395 0.555 2.395 0.39 1.605 0.39 1.605 0.33 2.455 0.33 2.455 0.495 3.27 0.495 3.27 0.435 3.33 0.435 ;
      POLYGON 3.01 1.13 2.97 1.13 2.97 1.305 2.525 1.305 2.525 1.225 2.89 1.225 2.89 1.05 3.01 1.05 ;
      POLYGON 2.79 1.125 2.26 1.125 2.26 1.38 1.495 1.38 1.495 1.16 1.7 1.16 1.7 0.715 1.165 0.715 1.165 0.78 1.105 0.78 1.105 0.655 1.7 0.655 1.7 0.49 1.76 0.49 1.76 1.22 1.555 1.22 1.555 1.32 2.2 1.32 2.2 1.065 2.73 1.065 2.73 0.915 2.79 0.915 ;
      POLYGON 0.76 1.02 0.68 1.02 0.68 0.815 0.425 0.815 0.425 0.735 0.68 0.735 0.68 0.54 0.76 0.54 ;
  END
END TLATSRXL

MACRO TLATX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATX1 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.708575 LAYER Metal1 ;
    ANTENNADIFFAREA 1.871125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.16875 LAYER Metal1 ;
      ANTENNAMAXAREACAR 10.124889 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 78.2755555 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.165 1.325 3.07 1.325 3.07 0.705 3.035 0.705 3.035 0.625 3.045 0.625 3.045 0.54 3.165 0.54 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.653475 LAYER Metal1 ;
    ANTENNADIFFAREA 1.871125 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.16875 LAYER Metal1 ;
      ANTENNAMAXAREACAR 9.79837025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 76.57777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.34 1.415 2.28 1.415 2.28 0.73 2.26 0.73 2.26 0.6 2.28 0.6 2.28 0.54 2.34 0.54 ;
    END
  END QN
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.78 1.94 1.28 ;
    END
  END G
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.635 1.025 0.46 1.025 0.46 0.62 0.54 0.62 0.54 0.725 0.635 0.725 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 1.77 0 1.77 0 1.65 0.375 1.65 0.375 1.285 0.435 1.285 0.435 1.65 1.235 1.65 1.235 1.54 1.355 1.54 1.355 1.65 2.075 1.65 2.075 1.295 2.135 1.295 2.135 1.65 2.84 1.65 2.84 0.965 2.9 0.965 2.9 1.65 3.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 0.06 2.9 0.06 2.9 0.52 2.84 0.52 2.84 0.06 2.105 0.06 2.105 0.52 2.045 0.52 2.045 0.06 1.38 0.06 1.38 0.2 1.32 0.2 1.32 0.06 0.52 0.06 0.52 0.2 0.46 0.2 0.46 0.06 0 0.06 0 -0.06 3.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.97 0.865 2.695 0.865 2.695 1.325 2.635 1.325 2.635 0.54 2.695 0.54 2.695 0.805 2.97 0.805 ;
      POLYGON 2.16 0.82 2.1 0.82 2.1 0.68 1.7 0.68 1.7 0.965 1.59 0.965 1.59 1.28 1.47 1.28 1.47 1.22 1.53 1.22 1.53 0.965 1.235 0.965 1.235 0.905 1.64 0.905 1.64 0.425 1.7 0.425 1.7 0.62 2.16 0.62 ;
      POLYGON 1.9 0.52 1.84 0.52 1.84 0.325 1.54 0.325 1.54 0.36 1.23 0.36 1.23 0.355 0.955 0.355 0.955 0.98 0.795 0.98 0.795 1.41 1.075 1.41 1.075 1.38 1.7 1.38 1.7 1.12 1.76 1.12 1.76 1.44 1.135 1.44 1.135 1.47 0.735 1.47 0.735 1.185 0.3 1.185 0.3 1.02 0.36 1.02 0.36 1.125 0.735 1.125 0.735 0.92 0.895 0.92 0.895 0.295 1.1 0.295 1.1 0.26 1.22 0.26 1.22 0.295 1.265 0.295 1.265 0.3 1.48 0.3 1.48 0.265 1.9 0.265 ;
      POLYGON 1.515 0.71 1.115 0.71 1.115 1.25 0.955 1.25 0.955 1.31 0.895 1.31 0.895 1.19 1.055 1.19 1.055 0.455 1.175 0.455 1.175 0.515 1.115 0.515 1.115 0.65 1.515 0.65 ;
      POLYGON 0.795 0.705 0.735 0.705 0.735 0.52 0.2 0.52 0.2 1.31 0.14 1.31 0.14 0.4 0.285 0.4 0.285 0.46 0.795 0.46 ;
  END
END TLATX1

MACRO TLATX2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATX2 0 0 ;
  SIZE 3.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 0.06 3.525 0.06 3.525 0.44 3.465 0.44 3.465 0.06 2.935 0.06 2.935 0.44 2.875 0.44 2.875 0.06 2.525 0.06 2.525 0.44 2.465 0.44 2.465 0.06 2.05 0.06 2.05 0.2 1.99 0.2 1.99 0.06 1.365 0.06 1.365 0.2 1.305 0.2 1.305 0.06 0.45 0.06 0.45 0.17 0.33 0.17 0.33 0.06 0 0.06 0 -0.06 3.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.6 1.77 0 1.77 0 1.65 0.33 1.65 0.33 1.345 0.39 1.345 0.39 1.65 1.33 1.65 1.33 1.375 1.45 1.375 1.45 1.435 1.39 1.435 1.39 1.65 2.055 1.65 2.055 1.185 2.115 1.185 2.115 1.65 2.465 1.65 2.465 0.915 2.525 0.915 2.525 1.65 2.875 1.65 2.875 0.915 2.935 0.915 2.935 1.65 3.465 1.65 3.465 0.915 3.525 0.915 3.525 1.65 3.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.59 0.815 0.565 0.815 0.565 1.085 0.36 1.085 0.36 0.735 0.59 0.735 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.835 0.815 2.015 1.085 ;
    END
  END G
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8628 LAYER Metal1 ;
    ANTENNADIFFAREA 2.35205 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.263475 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.0701205 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 55.8212355 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.34 0.54 2.32 0.54 2.32 1.305 2.26 1.305 2.26 0.41 2.34 0.41 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.9191 LAYER Metal1 ;
    ANTENNADIFFAREA 2.35205 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.263475 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.283803 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 56.93139775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.26 0.46 3.34 1.305 ;
    END
  END Q
  OBS
    LAYER Metal1 ;
      POLYGON 3.16 0.71 2.73 0.71 2.73 1.305 2.67 1.305 2.67 0.46 2.73 0.46 2.73 0.65 3.16 0.65 ;
      POLYGON 2.16 0.715 1.685 0.715 1.685 1.08 1.19 1.08 1.19 1.02 1.625 1.02 1.625 0.54 1.685 0.54 1.685 0.655 2.16 0.655 ;
      POLYGON 1.94 1.275 1.23 1.275 1.23 1.5 0.745 1.5 0.745 1.245 0.2 1.245 0.2 1.08 0.26 1.08 0.26 1.185 0.745 1.185 0.745 1 0.85 1 0.85 0.3 1.085 0.3 1.085 0.25 1.205 0.25 1.205 0.3 1.885 0.3 1.885 0.555 1.825 0.555 1.825 0.36 0.91 0.36 0.91 1.06 0.805 1.06 0.805 1.44 1.17 1.44 1.17 1.215 1.94 1.215 ;
      POLYGON 1.525 0.79 1.07 0.79 1.07 1.34 0.905 1.34 0.905 1.28 1.01 1.28 1.01 0.57 1.13 0.57 1.13 0.63 1.07 0.63 1.07 0.73 1.525 0.73 ;
      POLYGON 0.75 0.82 0.69 0.82 0.69 0.635 0.1 0.635 0.1 1.345 0.185 1.345 0.185 1.465 0.125 1.465 0.125 1.405 0.04 1.405 0.04 0.575 0.125 0.575 0.125 0.515 0.185 0.515 0.185 0.575 0.75 0.575 ;
  END
END TLATX2

MACRO TLATX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATX4 0 0 ;
  SIZE 4.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6486 LAYER Metal1 ;
    ANTENNADIFFAREA 3.4662 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.46215 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.73103975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 44.38169425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.95 0.585 2.48 0.585 2.48 1.025 2.77 1.025 2.77 1.355 2.71 1.355 2.71 1.085 2.36 1.085 2.36 1.355 2.26 1.355 2.26 0.98 2.42 0.98 2.42 0.465 2.48 0.465 2.48 0.525 2.89 0.525 2.89 0.465 2.95 0.465 ;
    END
  END QN
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6486 LAYER Metal1 ;
    ANTENNADIFFAREA 3.4662 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.46215 LAYER Metal1 ;
      ANTENNAMAXAREACAR 5.73103975 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 44.38169425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.13 1.355 1.07 1.355 1.07 1.025 0.72 1.025 0.72 1.355 0.66 1.355 0.66 0.79 0.68 0.79 0.68 0.585 0.54 0.585 0.54 0.465 0.6 0.465 0.6 0.525 1.01 0.525 1.01 0.465 1.07 0.465 1.07 0.585 0.74 0.585 0.74 0.965 1.13 0.965 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.54 1.065 4.46 1.065 4.46 0.92 4.235 0.92 4.235 0.79 4.54 0.79 ;
    END
  END D
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.26 0.46 0.34 0.96 ;
    END
  END G
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 1.77 0 1.77 0 1.65 0.455 1.65 0.455 0.965 0.515 0.965 0.515 1.65 0.865 1.65 0.865 1.125 0.925 1.125 0.925 1.65 1.275 1.65 1.275 0.965 1.335 0.965 1.335 1.65 1.685 1.65 1.685 1.125 1.745 1.125 1.745 1.65 2.095 1.65 2.095 0.965 2.155 0.965 2.155 1.65 2.505 1.65 2.505 1.185 2.565 1.185 2.565 1.65 2.915 1.65 2.915 0.965 2.975 0.965 2.975 1.65 3.355 1.65 3.355 1.165 3.415 1.165 3.415 1.65 4.31 1.65 4.31 1.165 4.37 1.165 4.37 1.65 4.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.8 0.06 4.4 0.06 4.4 0.2 4.34 0.2 4.34 0.06 3.74 0.06 3.74 0.2 3.68 0.2 3.68 0.06 3.215 0.06 3.215 0.17 3.095 0.17 3.095 0.06 2.745 0.06 2.745 0.17 2.625 0.17 2.625 0.06 2.275 0.06 2.275 0.17 2.155 0.17 2.155 0.06 1.805 0.06 1.805 0.17 1.685 0.17 1.685 0.06 1.335 0.06 1.335 0.17 1.215 0.17 1.215 0.06 0.865 0.06 0.865 0.17 0.745 0.17 0.745 0.06 0.28 0.06 0.28 0.2 0.22 0.2 0.22 0.06 0 0.06 0 -0.06 4.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.76 0.555 4.7 0.555 4.7 1.19 4.64 1.19 4.64 0.69 4.135 0.69 4.135 0.755 3.87 0.755 3.87 0.99 3.81 0.99 3.81 0.695 4.075 0.695 4.075 0.63 4.64 0.63 4.64 0.495 4.76 0.495 ;
      POLYGON 4.62 0.36 4.56 0.36 4.56 0.37 3.52 0.37 3.52 0.36 0.16 0.36 0.16 1.06 0.28 1.06 0.28 1.18 0.22 1.18 0.22 1.12 0.1 1.12 0.1 0.3 3.58 0.3 3.58 0.31 4.5 0.31 4.5 0.3 4.62 0.3 ;
      POLYGON 4.09 0.53 3.975 0.53 3.975 0.595 3.71 0.595 3.71 1.1 3.895 1.1 3.895 1.16 3.65 1.16 3.65 1.035 3.31 1.035 3.31 0.885 3.37 0.885 3.37 0.975 3.65 0.975 3.65 0.535 3.915 0.535 3.915 0.47 4.09 0.47 ;
      POLYGON 3.55 0.875 3.49 0.875 3.49 0.785 3.21 0.785 3.21 1.355 3.15 1.355 3.15 0.785 2.795 0.785 2.795 0.725 3.36 0.725 3.36 0.465 3.42 0.465 3.42 0.725 3.55 0.725 ;
      POLYGON 2.01 0.585 1.54 0.585 1.54 0.965 1.95 0.965 1.95 1.355 1.89 1.355 1.89 1.025 1.54 1.025 1.54 1.355 1.48 1.355 1.48 0.745 1.045 0.745 1.045 0.685 1.48 0.685 1.48 0.465 1.54 0.465 1.54 0.525 1.95 0.525 1.95 0.465 2.01 0.465 ;
  END
END TLATX4

MACRO TLATXL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TLATXL 0 0 ;
  SIZE 3.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.63505 LAYER Metal1 ;
    ANTENNADIFFAREA 1.65745 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1296 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.6161265 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 97.68518525 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 3.06 0.475 3.14 1.045 ;
    END
  END Q
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.68065 LAYER Metal1 ;
    ANTENNADIFFAREA 1.65745 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1296 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.9679785 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 99.18981475 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.35 1.49 2.155 1.49 2.155 1.36 2.27 1.36 2.27 0.405 2.35 0.405 ;
    END
  END QN
  PIN G
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 1.86 0.76 1.94 1.26 ;
    END
  END G
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.64 1.025 0.46 1.025 0.46 0.79 0.56 0.79 0.56 0.625 0.64 0.625 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 1.77 0 1.77 0 1.65 0.375 1.65 0.375 1.285 0.435 1.285 0.435 1.65 1.24 1.65 1.24 1.54 1.36 1.54 1.36 1.65 1.945 1.65 1.945 1.36 2.005 1.36 2.005 1.65 2.785 1.65 2.785 1.02 2.845 1.02 2.845 1.65 3.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.2 0.06 2.89 0.06 2.89 0.57 2.83 0.57 2.83 0.06 2.11 0.06 2.11 0.5 2.05 0.5 2.05 0.06 1.385 0.06 1.385 0.2 1.325 0.2 1.325 0.06 0.465 0.06 0.465 0.2 0.405 0.2 0.405 0.06 0 0.06 0 -0.06 3.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.915 0.855 2.685 0.855 2.685 0.985 2.64 0.985 2.64 1.045 2.58 1.045 2.58 0.925 2.625 0.925 2.625 0.475 2.685 0.475 2.685 0.795 2.915 0.795 ;
      POLYGON 2.17 0.685 2.05 0.685 2.05 0.66 1.705 0.66 1.705 0.97 1.6 0.97 1.6 1.28 1.48 1.28 1.48 1.22 1.54 1.22 1.54 0.97 1.24 0.97 1.24 0.91 1.645 0.91 1.645 0.43 1.705 0.43 1.705 0.6 2.17 0.6 ;
      POLYGON 1.905 0.5 1.845 0.5 1.845 0.33 1.545 0.33 1.545 0.36 0.96 0.36 0.96 0.98 0.8 0.98 0.8 1.41 1.06 1.41 1.06 1.38 1.71 1.38 1.71 1.32 1.77 1.32 1.77 1.44 1.12 1.44 1.12 1.47 0.74 1.47 0.74 1.185 0.3 1.185 0.3 1.02 0.36 1.02 0.36 1.125 0.74 1.125 0.74 0.92 0.9 0.92 0.9 0.3 1.105 0.3 1.105 0.265 1.225 0.265 1.225 0.3 1.485 0.3 1.485 0.27 1.905 0.27 ;
      POLYGON 1.525 0.69 1.12 0.69 1.12 1.25 0.96 1.25 0.96 1.31 0.9 1.31 0.9 1.19 1.06 1.19 1.06 0.46 1.18 0.46 1.18 0.52 1.12 0.52 1.12 0.63 1.525 0.63 ;
      POLYGON 0.8 0.71 0.74 0.71 0.74 0.525 0.2 0.525 0.2 1.31 0.14 1.31 0.14 0.405 0.23 0.405 0.23 0.465 0.8 0.465 ;
  END
END TLATXL

MACRO XNOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X1 0 0 ;
  SIZE 1.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.761425 LAYER Metal1 ;
    ANTENNADIFFAREA 0.831375 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06165 LAYER Metal1 ;
      ANTENNAMAXAREACAR 12.3507705 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 99.8540145 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.14 0.555 0.13 0.555 0.13 0.655 0.11 0.655 0.11 0.925 0.13 0.925 0.13 1.335 0.07 1.335 0.07 0.975 0.05 0.975 0.05 0.385 0.14 0.385 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.95370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.145 0.895 0.965 0.895 0.965 0.92 0.815 0.92 0.815 0.895 0.755 0.895 0.755 0.775 0.965 0.775 0.965 0.815 1.145 0.815 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.33333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.415 0.895 0.33 0.895 0.33 0.705 0.235 0.705 0.235 0.625 0.415 0.625 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 0.06 1.06 0.06 1.06 0.51 1 0.51 1 0.06 0.335 0.06 0.335 0.505 0.275 0.505 0.275 0.06 0 0.06 0 -0.06 1.4 -0.06 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.4 1.77 0 1.77 0 1.65 0.23 1.65 0.23 1.51 0.29 1.51 0.29 1.65 0.93 1.65 0.93 1.42 1.05 1.42 1.05 1.65 1.4 1.65 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 1.265 1.36 0.58 1.36 0.58 1.3 1.205 1.3 1.205 0.69 0.725 0.69 0.725 0.59 1.205 0.59 1.205 0.41 1.265 0.41 ;
      POLYGON 0.94 0.205 0.85 0.205 0.85 0.265 0.54 0.265 0.54 1.075 0.48 1.075 0.48 0.2 0.785 0.2 0.785 0.145 0.94 0.145 ;
      POLYGON 0.745 0.53 0.66 0.53 0.66 0.955 0.745 0.955 0.745 1.22 0.19 1.22 0.19 0.775 0.25 0.775 0.25 1.16 0.685 1.16 0.685 1.015 0.6 1.015 0.6 0.47 0.685 0.47 0.685 0.41 0.745 0.41 ;
  END
END XNOR2X1

MACRO XNOR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X2 0 0 ;
  SIZE 1.8 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.05355 LAYER Metal1 ;
    ANTENNADIFFAREA 1.0346 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0909 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.590209 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 91.980198 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.34 0.945 0.335 0.945 0.335 1.42 0.255 1.42 0.255 0.4 0.335 0.4 0.335 0.76 0.34 0.76 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.50925925 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.54 0.92 1.19 0.92 1.19 0.975 1.13 0.975 1.13 0.84 1.4 0.84 1.4 0.79 1.54 0.79 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.9444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.645 0.64 0.74 0.92 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.06 0.13 1.06 0.13 1.65 0.48 1.65 0.48 1.175 0.54 1.175 0.54 1.65 1.345 1.65 1.345 1.155 1.465 1.155 1.465 1.215 1.405 1.215 1.405 1.65 1.8 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.8 0.06 1.485 0.06 1.485 0.555 1.345 0.555 1.345 0.495 1.425 0.495 1.425 0.06 0.54 0.06 0.54 0.66 0.48 0.66 0.48 0.06 0.13 0.06 0.13 0.64 0.07 0.64 0.07 0.06 0 0.06 0 -0.06 1.8 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.69 1.15 1.58 1.15 1.58 1.095 1.245 1.095 1.245 1.44 0.885 1.44 0.885 1.38 1.185 1.38 1.185 1.035 1.58 1.035 1.58 1.03 1.62 1.03 1.62 0.715 1.225 0.715 1.225 0.78 1.125 0.78 1.125 0.655 1.585 0.655 1.585 0.49 1.645 0.49 1.645 0.655 1.69 0.655 ;
      POLYGON 1.335 0.39 0.845 0.39 0.845 0.54 0.865 0.54 0.865 1.075 0.845 1.075 0.845 1.15 0.785 1.15 0.785 1.02 0.805 1.02 0.805 0.6 0.785 0.6 0.785 0.33 1.335 0.33 ;
      POLYGON 1.05 1.28 0.62 1.28 0.62 1.115 0.405 1.115 0.405 0.82 0.47 0.82 0.47 1.055 0.68 1.055 0.68 1.22 0.99 1.22 0.99 0.49 1.05 0.49 ;
  END
END XNOR2X2

MACRO XNOR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2X4 0 0 ;
  SIZE 2.2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.37765 LAYER Metal1 ;
    ANTENNADIFFAREA 1.48025 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.8498575 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 59.059829 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.785 0.405 0.66 0.405 0.66 0.52 0.355 0.52 0.355 0.6 0.365 0.6 0.365 0.73 0.355 0.73 0.355 0.98 0.745 0.98 0.745 1.465 0.685 1.465 0.685 1.045 0.335 1.045 0.335 1.465 0.275 1.465 0.275 0.73 0.235 0.73 0.235 0.6 0.275 0.6 0.275 0.295 0.335 0.295 0.335 0.46 0.6 0.46 0.6 0.305 0.785 0.305 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.50165025 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.94 0.925 1.86 0.925 1.86 0.835 1.25 0.835 1.25 0.65 1.31 0.65 1.31 0.775 1.7 0.775 1.7 0.755 1.94 0.755 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.9444445 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.055 0.78 0.95 0.78 0.95 0.73 0.86 0.73 0.86 0.6 1.055 0.6 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.075 0.13 1.075 0.13 1.65 0.48 1.65 0.48 1.105 0.54 1.105 0.54 1.65 0.89 1.65 0.89 1.225 0.95 1.225 0.95 1.65 1.795 1.65 1.795 1.105 1.855 1.105 1.855 1.65 2.2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.2 0.06 1.81 0.06 1.81 0.515 1.69 0.515 1.69 0.06 0.95 0.06 0.95 0.405 0.845 0.405 0.845 0.06 0.54 0.06 0.54 0.4 0.44 0.4 0.44 0.06 0.13 0.06 0.13 0.515 0.07 0.515 0.07 0.06 0 0.06 0 -0.06 2.2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.09 1.195 2.03 1.195 2.03 0.665 1.39 0.665 1.39 0.605 1.955 0.605 1.955 0.405 2.09 0.405 ;
      POLYGON 1.79 1.035 1.695 1.035 1.695 1.005 1.37 1.005 1.37 1.165 1.25 1.165 1.25 1.01 1.13 1.01 1.13 0.41 1.19 0.41 1.19 0.945 1.695 0.945 1.695 0.915 1.79 0.915 ;
      POLYGON 1.545 1.405 1.09 1.405 1.09 1.165 0.805 1.165 0.805 0.92 0.615 0.92 0.615 0.605 0.72 0.605 0.72 0.465 1.01 0.465 1.01 0.23 1.415 0.23 1.415 0.515 1.355 0.515 1.355 0.29 1.07 0.29 1.07 0.525 0.78 0.525 0.78 0.665 0.68 0.665 0.68 0.86 0.865 0.86 0.865 1.105 1.15 1.105 1.15 1.345 1.485 1.345 1.485 1.12 1.545 1.12 ;
  END
END XNOR2X4

MACRO XNOR2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2XL 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.825575 LAYER Metal1 ;
    ANTENNADIFFAREA 0.85685 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.98714 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 137.16049375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.195 0.705 0.15 0.705 0.15 1.11 0.09 1.11 0.09 0.73 0.06 0.73 0.06 0.6 0.135 0.6 0.135 0.485 0.195 0.485 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 5.04629625 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.315 0.935 0.89 0.935 0.89 0.855 1.03 0.855 1.03 0.815 1.315 0.815 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.4074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 0.92 0.395 0.92 0.395 0.665 0.475 0.665 0.475 0.79 0.54 0.79 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.37 1.65 0.37 1.38 0.43 1.38 0.43 1.65 1.095 1.65 1.095 1.405 1.215 1.405 1.215 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.275 0.06 1.275 0.55 1.14 0.55 1.14 0.49 1.215 0.49 1.215 0.06 0.4 0.06 0.4 0.58 0.34 0.58 0.34 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.435 1.11 1.02 1.11 1.02 1.45 0.65 1.45 0.65 1.39 0.96 1.39 0.96 1.05 1.375 1.05 1.375 0.715 0.95 0.715 0.95 0.775 0.89 0.775 0.89 0.655 1.375 0.655 1.375 0.485 1.435 0.485 ;
      POLYGON 1.115 0.385 0.605 0.385 0.605 0.635 0.66 0.635 0.66 1.07 0.605 1.07 0.605 1.17 0.545 1.17 0.545 1.01 0.6 1.01 0.6 0.7 0.545 0.7 0.545 0.325 1.115 0.325 ;
      POLYGON 0.815 1.31 0.21 1.31 0.21 0.81 0.27 0.81 0.27 1.25 0.755 1.25 0.755 0.485 0.815 0.485 ;
  END
END XNOR2XL

MACRO XNOR3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR3X1 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 4.065 0.06 4.065 0.64 4.005 0.64 4.005 0.06 1.04 0.06 1.04 0.17 0.92 0.17 0.92 0.135 0.425 0.135 0.425 0.17 0.305 0.17 0.305 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.335 1.65 0.335 1.365 0.395 1.365 0.395 1.65 1.025 1.65 1.025 1.54 1.145 1.54 1.145 1.575 4.005 1.575 4.005 1.01 4.065 1.01 4.065 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.045 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.73333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.365 0.935 3.235 0.935 3.235 0.725 2.925 0.725 2.925 0.665 3.295 0.665 3.295 0.815 3.365 0.815 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.071775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.4242425 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 1.055 0.46 1.055 0.46 0.75 0.41 0.75 0.41 0.605 0.49 0.605 0.49 0.67 0.54 0.67 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.026775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.4985995 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.105 0.07 1.105 0.07 0.92 0.06 0.92 0.06 0.79 0.07 0.79 0.07 0.615 0.15 0.615 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.723625 LAYER Metal1 ;
    ANTENNADIFFAREA 2.94 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.121725 LAYER Metal1 ;
      ANTENNAMAXAREACAR 22.375231 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 158.15157125 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.365 0.99 4.24 0.99 4.24 0.93 4.305 0.93 4.305 0.515 4.235 0.515 4.235 0.435 4.365 0.435 ;
    END
  END Y
  OBS
    LAYER Metal1 ;
      POLYGON 4.16 0.86 3.905 0.86 3.905 1.29 3.17 1.29 3.17 1.23 3.845 1.23 3.845 0.47 3.14 0.47 3.14 0.41 3.905 0.41 3.905 0.8 4.1 0.8 4.1 0.74 4.16 0.74 ;
      POLYGON 3.745 0.65 3.705 0.65 3.705 1.02 3.745 1.02 3.745 1.1 3.625 1.1 3.625 0.57 3.745 0.57 ;
      POLYGON 3.525 1.13 2.01 1.13 2.01 1.07 2.485 1.07 2.485 0.45 2.2 0.45 2.2 0.39 2.545 0.39 2.545 1.07 3.465 1.07 3.465 0.63 3.405 0.63 3.405 0.57 3.525 0.57 ;
      POLYGON 3.055 0.97 2.765 0.97 2.765 0.48 2.995 0.48 2.995 0.54 2.825 0.54 2.825 0.91 3.055 0.91 ;
      RECT 1.585 1.23 3.055 1.29 ;
      RECT 1.185 0.23 2.715 0.29 ;
      RECT 1.29 1.39 2.715 1.45 ;
      POLYGON 2.385 0.705 2.09 0.705 2.09 0.83 2.01 0.83 2.01 0.625 2.385 0.625 ;
      POLYGON 2.015 0.45 1.91 0.45 1.91 1.13 0.955 1.13 0.955 1.395 0.495 1.395 0.495 1.265 0.16 1.265 0.16 1.325 0.1 1.325 0.1 1.205 0.25 1.205 0.25 0.515 0.07 0.515 0.07 0.295 0.76 0.295 0.76 0.235 0.82 0.235 0.82 0.355 0.13 0.355 0.13 0.455 0.31 0.455 0.31 1.205 0.555 1.205 0.555 1.335 0.895 1.335 0.895 1.07 1.85 1.07 1.85 0.39 2.015 0.39 ;
      POLYGON 1.75 0.65 1.67 0.65 1.67 0.63 1.57 0.63 1.57 0.81 1.385 0.81 1.385 0.73 1.49 0.73 1.49 0.55 1.67 0.55 1.67 0.53 1.75 0.53 ;
      POLYGON 1.675 0.97 1.225 0.97 1.225 0.39 1.57 0.39 1.57 0.45 1.285 0.45 1.285 0.91 1.675 0.91 ;
      POLYGON 0.87 0.885 0.735 0.885 0.735 1.155 0.775 1.155 0.775 1.235 0.655 1.235 0.655 0.535 0.57 0.535 0.57 0.455 0.735 0.455 0.735 0.805 0.87 0.805 ;
  END
END XNOR3X1

MACRO XNOR3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR3XL 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.35 1.65 0.35 1.36 0.41 1.36 0.41 1.65 1.02 1.65 1.02 1.54 1.14 1.54 1.14 1.65 4.005 1.65 4.005 1.025 4.065 1.025 4.065 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.469775 LAYER Metal1 ;
    ANTENNADIFFAREA 2.89955 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.109125 LAYER Metal1 ;
      ANTENNAMAXAREACAR 22.6325315 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 176.65979375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.365 1.1 4.24 1.1 4.24 1.04 4.305 1.04 4.305 0.705 4.235 0.705 4.235 0.625 4.24 0.625 4.24 0.57 4.365 0.57 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.023175 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.5080905 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.175 1.1 0.095 1.1 0.095 0.92 0.06 0.92 0.06 0.79 0.095 0.79 0.095 0.635 0.175 0.635 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0675 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 2.57777775 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.54 1.1 0.46 1.1 0.46 0.78 0.435 0.78 0.435 0.625 0.515 0.625 0.515 0.7 0.54 0.7 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.045 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.73333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.365 0.935 3.035 0.935 3.035 0.725 2.925 0.725 2.925 0.665 3.095 0.665 3.095 0.815 3.165 0.815 3.165 0.875 3.365 0.875 ;
    END
  END C
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 4.065 0.06 4.065 0.66 4.005 0.66 4.005 0.06 1.065 0.06 1.065 0.17 0.945 0.17 0.945 0.06 0.44 0.06 0.44 0.17 0.32 0.17 0.32 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 4.16 0.925 3.905 0.925 3.905 1.29 3.17 1.29 3.17 1.23 3.845 1.23 3.845 0.47 3.14 0.47 3.14 0.41 3.905 0.41 3.905 0.865 4.1 0.865 4.1 0.805 4.16 0.805 ;
      POLYGON 3.745 0.65 3.705 0.65 3.705 1.02 3.745 1.02 3.745 1.1 3.625 1.1 3.625 0.57 3.745 0.57 ;
      POLYGON 3.525 1.13 2.035 1.13 2.035 1.07 2.51 1.07 2.51 0.465 2.225 0.465 2.225 0.405 2.57 0.405 2.57 1.07 3.465 1.07 3.465 0.63 3.405 0.63 3.405 0.57 3.525 0.57 ;
      POLYGON 2.995 0.54 2.825 0.54 2.825 0.91 2.935 0.91 2.935 0.97 2.765 0.97 2.765 0.48 2.995 0.48 ;
      RECT 1.58 1.23 2.935 1.29 ;
      RECT 1.21 0.23 2.74 0.29 ;
      RECT 1.285 1.39 2.74 1.45 ;
      POLYGON 2.41 0.685 2.115 0.685 2.115 0.81 2.035 0.81 2.035 0.605 2.41 0.605 ;
      POLYGON 2.04 0.45 1.935 0.45 1.935 1.13 0.95 1.13 0.95 1.44 0.51 1.44 0.51 1.26 0.175 1.26 0.175 1.32 0.115 1.32 0.115 1.2 0.275 1.2 0.275 0.535 0.085 0.535 0.085 0.315 0.785 0.315 0.785 0.255 0.845 0.255 0.845 0.375 0.145 0.375 0.145 0.475 0.335 0.475 0.335 1.2 0.57 1.2 0.57 1.38 0.89 1.38 0.89 1.07 1.875 1.07 1.875 0.39 2.04 0.39 ;
      POLYGON 1.775 0.64 1.695 0.64 1.695 0.63 1.595 0.63 1.595 0.81 1.38 0.81 1.38 0.73 1.515 0.73 1.515 0.55 1.695 0.55 1.695 0.52 1.775 0.52 ;
      POLYGON 1.67 0.97 1.22 0.97 1.22 0.39 1.595 0.39 1.595 0.45 1.28 0.45 1.28 0.91 1.67 0.91 ;
      POLYGON 0.865 0.885 0.75 0.885 0.75 1.2 0.79 1.2 0.79 1.28 0.67 1.28 0.67 0.555 0.595 0.555 0.595 0.475 0.75 0.475 0.75 0.805 0.865 0.805 ;
  END
END XNOR3XL

MACRO XOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X1 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.822225 LAYER Metal1 ;
    ANTENNADIFFAREA 0.91115 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.06165 LAYER Metal1 ;
      ANTENNAMAXAREACAR 13.336983 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 107.83455 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.2 1.29 0.14 1.29 0.14 1.11 0.06 1.11 0.06 0.98 0.14 0.98 0.14 0.38 0.2 0.38 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.14814825 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.405 0.87 1.165 0.87 1.165 0.92 1.035 0.92 1.035 0.87 0.67 0.87 0.67 0.775 1.405 0.775 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 11.0185185 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.565 0.54 0.49 0.54 0.49 0.85 0.41 0.85 0.41 0.41 0.565 0.41 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.345 1.65 0.345 1.49 0.465 1.49 0.465 1.65 1.165 1.65 1.165 1.17 1.225 1.17 1.225 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.245 0.06 1.245 0.55 1.185 0.55 1.185 0.06 0.465 0.06 0.465 0.215 0.345 0.215 0.345 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.525 1.01 1.43 1.01 1.43 1.195 1.37 1.195 1.37 1.11 0.89 1.11 0.89 1.005 0.815 1.005 0.815 0.945 0.95 0.945 0.95 1.05 1.37 1.05 1.37 0.945 1.465 0.945 1.465 0.575 1.39 0.575 1.39 0.455 1.45 0.455 1.45 0.515 1.525 0.515 ;
      POLYGON 1.245 0.715 0.61 0.715 0.61 1.135 0.62 1.135 0.62 1.27 0.55 1.27 0.55 0.655 0.66 0.655 0.66 0.455 0.73 0.455 0.73 0.655 1.245 0.655 ;
      POLYGON 0.935 0.55 0.875 0.55 0.875 0.335 0.33 0.335 0.33 1.33 0.765 1.33 0.765 1.14 0.825 1.14 0.825 1.39 0.27 1.39 0.27 0.275 0.935 0.275 ;
  END
END XOR2X1

MACRO XOR2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X2 0 0 ;
  SIZE 2 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.0182 LAYER Metal1 ;
    ANTENNADIFFAREA 1.164775 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0909 LAYER Metal1 ;
      ANTENNAMAXAREACAR 11.20132025 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 91.320132 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.435 0.555 0.34 0.555 0.34 1.155 0.435 1.155 0.435 1.275 0.375 1.275 0.375 1.215 0.28 1.215 0.28 0.73 0.26 0.73 0.26 0.6 0.28 0.6 0.28 0.495 0.375 0.495 0.375 0.435 0.435 0.435 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.45370375 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.785 0.875 1.565 0.875 1.565 0.895 1.435 0.895 1.435 0.885 1.06 0.885 1.06 0.825 1.335 0.825 1.335 0.815 1.785 0.815 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.8 1.195 0.72 1.195 0.72 0.895 0.6 0.895 0.6 0.815 0.8 0.815 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 1.77 0 1.77 0 1.65 0.12 1.65 0.12 0.985 0.18 0.985 0.18 1.65 0.58 1.65 0.58 1.54 0.7 1.54 0.7 1.65 1.52 1.65 1.52 1.17 1.58 1.17 1.58 1.65 2 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2 0.06 1.625 0.06 1.625 0.55 1.565 0.55 1.565 0.06 0.64 0.06 0.64 0.52 0.58 0.52 0.58 0.06 0.18 0.06 0.18 0.52 0.12 0.52 0.12 0.06 0 0.06 0 -0.06 2 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.945 1.07 1.785 1.07 1.785 1.195 1.725 1.195 1.725 1.07 1.42 1.07 1.42 1.42 1.22 1.42 1.22 1.36 1.36 1.36 1.36 1.01 1.885 1.01 1.885 0.575 1.77 0.575 1.77 0.455 1.83 0.455 1.83 0.515 1.945 0.515 ;
      POLYGON 1.625 0.715 0.96 0.715 0.96 1.195 0.9 1.195 0.9 0.485 1.02 0.485 1.02 0.545 0.96 0.545 0.96 0.655 1.625 0.655 ;
      POLYGON 1.315 0.55 1.255 0.55 1.255 0.385 0.8 0.385 0.8 0.715 0.5 0.715 0.5 0.995 0.62 0.995 0.62 1.295 1.06 1.295 1.06 1.2 1.165 1.2 1.165 1.14 1.225 1.14 1.225 1.26 1.12 1.26 1.12 1.355 0.56 1.355 0.56 1.055 0.44 1.055 0.44 0.655 0.74 0.655 0.74 0.325 1.315 0.325 ;
  END
END XOR2X2

MACRO XOR2X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2X4 0 0 ;
  SIZE 2.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.3541 LAYER Metal1 ;
    ANTENNADIFFAREA 1.614025 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.1755 LAYER Metal1 ;
      ANTENNAMAXAREACAR 7.7156695 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 61.880342 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.745 0.45 0.7 0.45 0.7 0.61 0.32 0.61 0.32 0.98 0.34 0.98 0.34 1.075 0.7 1.075 0.7 1.345 0.745 1.345 0.745 1.465 0.685 1.465 0.685 1.405 0.64 1.405 0.64 1.135 0.335 1.135 0.335 1.465 0.26 1.465 0.26 0.56 0.245 0.56 0.245 0.5 0.365 0.5 0.365 0.55 0.64 0.55 0.64 0.39 0.685 0.39 0.685 0.33 0.745 0.33 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.04545 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 3.82838275 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.205 0.745 2.125 0.745 2.125 0.705 1.745 0.705 1.745 0.625 2.205 0.625 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 10.74074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        RECT 0.96 0.71 1.165 1.085 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 1.77 0 1.77 0 1.65 0.07 1.65 0.07 1.075 0.13 1.075 0.13 1.65 0.48 1.65 0.48 1.235 0.54 1.235 0.54 1.65 0.86 1.65 0.86 1.375 0.98 1.375 0.98 1.435 0.92 1.435 0.92 1.65 2.02 1.65 2.02 1.125 2.08 1.125 2.08 1.65 2.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 2.4 0.06 2.05 0.06 2.05 0.305 2.11 0.305 2.11 0.365 1.99 0.365 1.99 0.06 0.95 0.06 0.95 0.45 0.89 0.45 0.89 0.06 0.54 0.06 0.54 0.45 0.48 0.45 0.48 0.06 0.13 0.06 0.13 0.45 0.07 0.45 0.07 0.06 0 0.06 0 -0.06 2.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 2.365 0.905 2.285 0.905 2.285 1.15 2.225 1.15 2.225 0.845 2.305 0.845 2.305 0.525 1.645 0.525 1.645 0.805 1.825 0.805 1.825 0.865 1.585 0.865 1.585 0.665 1.485 0.665 1.485 0.725 1.425 0.725 1.425 0.605 1.585 0.605 1.585 0.465 2.225 0.465 2.225 0.3 2.285 0.3 2.285 0.465 2.365 0.465 ;
      POLYGON 2.045 0.905 1.985 0.905 1.985 1.025 1.325 1.025 1.325 1.195 1.265 1.195 1.265 0.445 1.385 0.445 1.385 0.505 1.325 0.505 1.325 0.965 1.925 0.965 1.925 0.845 2.045 0.845 ;
      POLYGON 1.73 1.355 1.105 1.355 1.105 1.245 0.8 1.245 0.8 0.77 0.59 0.77 0.59 0.71 0.8 0.71 0.8 0.55 1.105 0.55 1.105 0.285 1.575 0.285 1.575 0.305 1.645 0.305 1.645 0.365 1.525 0.365 1.525 0.345 1.165 0.345 1.165 0.61 0.86 0.61 0.86 1.185 1.165 1.185 1.165 1.295 1.67 1.295 1.67 1.235 1.73 1.235 ;
  END
END XOR2X4

MACRO XOR2XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2XL 0 0 ;
  SIZE 1.6 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.8073 LAYER Metal1 ;
    ANTENNADIFFAREA 0.865 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0486 LAYER Metal1 ;
      ANTENNAMAXAREACAR 16.611111 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 136.85185175 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.15 1.18 0.07 1.18 0.07 0.735 0.06 0.735 0.06 0.59 0.07 0.59 0.07 0.44 0.15 0.44 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0324 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 8.24074075 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.37 0.895 0.765 0.895 0.765 1.025 0.705 1.025 0.705 0.8 1.37 0.8 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0162 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.611111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.565 0.54 0.45 0.54 0.45 0.95 0.37 0.95 0.37 0.41 0.565 0.41 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 1.77 0 1.77 0 1.65 0.325 1.65 0.325 1.465 0.385 1.465 0.385 1.65 1.15 1.65 1.15 1.155 1.21 1.155 1.21 1.65 1.6 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 1.6 0.06 1.31 0.06 1.31 0.535 1.25 0.535 1.25 0.06 0.355 0.06 0.355 0.225 0.295 0.225 0.295 0.06 0 0.06 0 -0.06 1.6 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  OBS
    LAYER Metal1 ;
      POLYGON 1.515 1.055 1.415 1.055 1.415 1.18 1.355 1.18 1.355 1.055 0.955 1.055 0.955 1.435 0.895 1.435 0.895 0.995 1.455 0.995 1.455 0.44 1.515 0.44 ;
      POLYGON 1.3 0.69 0.635 0.69 0.635 1.025 0.605 1.025 0.605 1.18 0.545 1.18 0.545 0.955 0.575 0.955 0.575 0.63 0.67 0.63 0.67 0.435 0.73 0.435 0.73 0.63 1.3 0.63 ;
      POLYGON 0.985 0.535 0.925 0.535 0.925 0.345 0.29 0.345 0.29 1.275 0.755 1.275 0.755 1.125 0.815 1.125 0.815 1.335 0.23 1.335 0.23 0.285 0.985 0.285 ;
  END
END XOR2XL

MACRO XOR3X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR3X1 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 4.065 0.06 4.065 0.66 4.005 0.66 4.005 0.06 1.14 0.06 1.14 0.17 1.02 0.17 1.02 0.135 0.425 0.135 0.425 0.17 0.305 0.17 0.305 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.045 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.73333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.365 0.935 3.235 0.935 3.235 0.725 2.925 0.725 2.925 0.665 3.295 0.665 3.295 0.815 3.365 0.815 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0868 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.071775 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.20933475 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 12.831766 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.64 0.895 0.43 0.895 0.43 0.525 0.51 0.525 0.51 0.815 0.64 0.815 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.026775 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 6.4985995 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.17 1.085 0.09 1.085 0.09 0.92 0.06 0.92 0.06 0.79 0.09 0.79 0.09 0.615 0.17 0.615 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.387225 LAYER Metal1 ;
    ANTENNADIFFAREA 2.95605 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.12105 LAYER Metal1 ;
      ANTENNAMAXAREACAR 19.720983 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 149.1697645 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.365 1.085 4.24 1.085 4.24 1.025 4.305 1.025 4.305 0.705 4.235 0.705 4.235 0.625 4.24 0.625 4.24 0.57 4.365 0.57 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.235 1.65 0.235 1.345 0.395 1.345 0.395 1.65 1.125 1.65 1.125 1.54 1.245 1.54 1.245 1.65 4.005 1.65 4.005 1.025 4.065 1.025 4.065 1.65 4.4 1.65 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VDD:%:VDD!]" ;
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.16 0.925 3.905 0.925 3.905 1.29 3.17 1.29 3.17 1.23 3.845 1.23 3.845 0.47 3.14 0.47 3.14 0.41 3.905 0.41 3.905 0.865 4.1 0.865 4.1 0.805 4.16 0.805 ;
      POLYGON 3.745 0.65 3.705 0.65 3.705 1.02 3.745 1.02 3.745 1.1 3.625 1.1 3.625 0.57 3.745 0.57 ;
      POLYGON 3.525 1.13 2.11 1.13 2.11 1.07 2.585 1.07 2.585 0.45 2.27 0.45 2.27 0.39 2.645 0.39 2.645 1.07 3.465 1.07 3.465 0.63 3.405 0.63 3.405 0.57 3.525 0.57 ;
      POLYGON 3.055 0.97 2.765 0.97 2.765 0.48 2.995 0.48 2.995 0.54 2.825 0.54 2.825 0.91 3.055 0.91 ;
      RECT 1.685 1.23 3.055 1.29 ;
      RECT 1.285 0.23 2.815 0.29 ;
      RECT 1.39 1.39 2.815 1.45 ;
      POLYGON 2.485 0.705 2.19 0.705 2.19 0.83 2.11 0.83 2.11 0.625 2.485 0.625 ;
      POLYGON 2.115 0.45 2.01 0.45 2.01 1.13 1.055 1.13 1.055 1.245 0.135 1.245 0.135 1.305 0.075 1.305 0.075 1.185 0.27 1.185 0.27 0.515 0.07 0.515 0.07 0.295 0.86 0.295 0.86 0.235 0.92 0.235 0.92 0.355 0.13 0.355 0.13 0.455 0.33 0.455 0.33 1.185 0.995 1.185 0.995 1.07 1.95 1.07 1.95 0.39 2.115 0.39 ;
      POLYGON 1.85 0.65 1.77 0.65 1.77 0.63 1.67 0.63 1.67 0.81 1.485 0.81 1.485 0.73 1.59 0.73 1.59 0.55 1.77 0.55 1.77 0.53 1.85 0.53 ;
      POLYGON 1.775 0.97 1.325 0.97 1.325 0.39 1.67 0.39 1.67 0.45 1.385 0.45 1.385 0.91 1.775 0.91 ;
      POLYGON 0.86 0.725 0.82 0.725 0.82 1.075 0.655 1.075 0.655 0.995 0.74 0.995 0.74 0.715 0.71 0.715 0.71 0.535 0.67 0.535 0.67 0.455 0.79 0.455 0.79 0.645 0.86 0.645 ;
  END
END XOR3X1

MACRO XOR3XL
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR3XL 0 0 ;
  SIZE 4.4 BY 1.71 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    NETEXPR "VSS VSS!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 0.06 4.065 0.06 4.065 0.66 4.005 0.66 4.005 0.06 1.065 0.06 1.065 0.17 0.945 0.17 0.945 0.06 0.44 0.06 0.44 0.17 0.32 0.17 0.32 0.06 0 0.06 0 -0.06 4.4 -0.06 ;
    END
    PROPERTY DB_Inherited_Net_Expr "[@VSS:%:VSS!]" ;
  END VSS
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.045 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 4.73333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 3.365 0.935 3.235 0.935 3.235 0.725 2.925 0.725 2.925 0.665 3.295 0.665 3.295 0.815 3.365 0.815 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.0892 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0675 LAYER Metal1 ;
      ANTENNAMAXAREACAR 1.3214815 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 13.911111 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.57 1.085 0.435 1.085 0.435 0.64 0.515 0.64 0.515 1.005 0.57 1.005 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.0225 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 7.73333325 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 0.175 1.115 0.095 1.115 0.095 0.92 0.06 0.92 0.06 0.79 0.095 0.79 0.095 0.65 0.175 0.65 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.3408 LAYER Metal1 ;
    ANTENNADIFFAREA 2.82975 LAYER Metal1 ;
    ANTENNAMODEL OXIDE1 ;
      ANTENNAGATEAREA 0.107775 LAYER Metal1 ;
      ANTENNAMAXAREACAR 21.71932275 LAYER Metal1 ;
      ANTENNAMAXSIDEAREACAR 170.4244955 LAYER Metal1 ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.365 1.1 4.24 1.1 4.24 1.04 4.305 1.04 4.305 0.705 4.235 0.705 4.235 0.625 4.24 0.625 4.24 0.57 4.365 0.57 ;
    END
  END Y
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    NETEXPR "VDD VDD!" ;
    PORT
      LAYER Metal1 ;
        POLYGON 4.4 1.77 0 1.77 0 1.65 0.35 1.65 0.35 1.375 0.41 1.375 0.41 1.65 1.02 1.65 1.02 1.54 1.14 1.54 1.14 1.65 4.005 1.65 4.005 1.025 4.065 1.025 4.065 1.65 4.4 1.65 ;
    END
  END VDD
  OBS
    LAYER Metal1 ;
      POLYGON 4.16 0.925 3.905 0.925 3.905 1.29 3.17 1.29 3.17 1.23 3.845 1.23 3.845 0.47 3.14 0.47 3.14 0.41 3.905 0.41 3.905 0.865 4.1 0.865 4.1 0.805 4.16 0.805 ;
      POLYGON 3.745 0.65 3.705 0.65 3.705 1.02 3.745 1.02 3.745 1.1 3.625 1.1 3.625 0.57 3.745 0.57 ;
      POLYGON 3.525 1.13 2.035 1.13 2.035 1.07 2.51 1.07 2.51 0.45 2.195 0.45 2.195 0.39 2.57 0.39 2.57 1.07 3.465 1.07 3.465 0.63 3.405 0.63 3.405 0.57 3.525 0.57 ;
      POLYGON 3.055 0.97 2.765 0.97 2.765 0.48 2.995 0.48 2.995 0.54 2.825 0.54 2.825 0.91 3.055 0.91 ;
      RECT 1.58 1.23 3.055 1.29 ;
      RECT 1.21 0.23 2.74 0.29 ;
      RECT 1.285 1.39 2.74 1.45 ;
      POLYGON 2.41 0.685 2.115 0.685 2.115 0.81 2.035 0.81 2.035 0.605 2.41 0.605 ;
      POLYGON 2.04 0.45 1.935 0.45 1.935 1.13 0.95 1.13 0.95 1.425 0.51 1.425 0.51 1.275 0.175 1.275 0.175 1.335 0.115 1.335 0.115 1.215 0.275 1.215 0.275 0.55 0.085 0.55 0.085 0.33 0.785 0.33 0.785 0.27 0.845 0.27 0.845 0.39 0.145 0.39 0.145 0.49 0.335 0.49 0.335 1.215 0.57 1.215 0.57 1.365 0.89 1.365 0.89 1.07 1.875 1.07 1.875 0.39 2.04 0.39 ;
      POLYGON 1.775 0.64 1.695 0.64 1.695 0.63 1.595 0.63 1.595 0.81 1.38 0.81 1.38 0.73 1.515 0.73 1.515 0.55 1.695 0.55 1.695 0.52 1.775 0.52 ;
      POLYGON 1.67 0.97 1.22 0.97 1.22 0.39 1.595 0.39 1.595 0.45 1.28 0.45 1.28 0.91 1.67 0.91 ;
      POLYGON 0.79 0.75 0.75 0.75 0.75 1.185 0.79 1.185 0.79 1.265 0.67 1.265 0.67 0.75 0.635 0.75 0.635 0.57 0.595 0.57 0.595 0.49 0.715 0.49 0.715 0.67 0.79 0.67 ;
  END
END XOR3XL

END LIBRARY
